��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b����K=&no��|�.�0����4�C�wI���V��ƨMU���GW��x[`O��+l��|@��������|�d%A���'�6%��gf9��1NSv���Hf��nc�_���ȿo�|DJs/ �~r]�����5��ʉb\�i�5��}��'j|��"/��<����"��o� �6Z�'O"�9�������$�CmOL��e��$��u��Ue�����.�����ȦԄ6S�W�FL�=-�]<�N�L�ǌ�����Z�=��2�%��j[\��zWm�I�ƫ�e/���zS�'NFP�'����+w�7���_-�_��o$^%�P�·�G���U:|*��xoo�&{m�u�͵m�{^��ڧW��7T������m�ye(ͮ1���W�F/���,]���K,���h[����G����/P`������Z���H���_�#?��S�v+#dP0�>���+�Q8����Aw`*;�fQ�;��B�Y?K(�K�/ ��pX���t�&z�,��GԺ�����=_3}s�����j���3�O�����5�����9P%J���ĉN���(|�-I�z��VdҎC"�B��kN�U����l�})Ч�\S�(!<#���	3"�@���[C��6_SbZ�Z�_=Ի�$51ES~j��l�@f1�NX62�E<��,�*g�5
��U��D�C^#��u�l�a�iY۸M�Ģ����x�e߮�["d�Q�,i3�q�=�Ǩ�:1�΂�12P���m¤�z�/K{�՞����H-{�� F�P�/3�u��1OP7���-��,U���
>i��� <�4� c=M+�5>g�n..�Uڥ%цsK|}�7nh��O��/����0ON��@B5@J�c)OF���w�D7W��Q��Xl��6n�ӥ�7�G�����Ս���(B�Mn/b�@�(��V�d2�\�^G���'i��w�~�sJg�7�A�$��q�ӌ6�t�KsRZ9n��P?E�M�e�֭��]ȯ�����E��I��Ig�,�G��V���"���,��1�n�a�p-��?��&cE�&��SH+x]Q�u��g�\�s|e}�6��|�h�g��Ŭb�+$N�=O���8�?��>�Q}ȽM4̅���G�T���@��?U�uyq9C��p�I>�cS9R�ط��J���J�k���JN9�/�/�]� ׀�G�U��4�C�H_���)d�>=
m��Ҿ{C�f�It��2�pt����5��P�K?6p��J�u�}"?��N������p�x���4)�� �A��f�t�bxL��,zQ�dB�b��������?`~�~�����$8'��G{����ǆ��u��j��Q�V����6�dЀ���5,Aa<�h�*/:��;�c�����`%���[�ӵ_�ɩyi����[�7-_��3��*+�q 6>o�����+m�e1��+�{I_n�ŵ�N�l%V�Hm{�z;�[�s1�d�������0��pɦ��������S07Jd)F�-�QGK.��{@ ~�RR;t���*��c���X����¡ÐIB�W�'���2�=s *3:���ѡ$8N�r�q�᳊�0<�����"W̞i�����8��"�{�;M
l�Nl���RX�2	���1�&��j/#X;��:Qr�slQy:v!۱3$A2�v�ߛ�OGS�^>�=J�S�	n�.eV,�+Θ?+��1�p��$�F�)K8��G�[�r��cmS�k�ԇA�&��	��,��J�Q�KژF��/6m0y����oO�ا;�j�#y7�=�N'J]��Xn���~ �C*Y��Nߏ!�"k����^05H������~�nF/���{x0��/4'��G%�XtO9	��M�$lQn�
�
���S�P>�g�O��N�$Jya="�0�t�O��Ӛ���qq3�w����Q�ђ���@/��Е��.0h&4,�'r�o�j�� h[6&�^�*�~>�Ί�9bZ�%�1]T�	(
�=vhmZ����Rt��Y�` ��&`�5��d���4p��!	t[��T���x�����ŕ�	}q�2�ByX}�9�U��(��o���3���q��#������Xf���<�}vCo�54Pq�4WT30������ŖA9�O�9�l�Fk�tɔ�N�M���s����9��$`U�5y5�8n�Gi��jEp��i�e46��4tٮ���y�'�8`O�x�0P�~��2j��T�{D=�B�~\/�OZd0"��)��ܾ	��Z<n�V��DU2���O+�0Mh�DX�<c�	�0��-X�D��/�v���]��������H��+/Jf�Q��qv5t�W_���\P�w�p$`3y(s��d����3�{jR���~j4	���GX����ǰ`��y�`�=��?8T	�#pL�l3��U��{�\�W�i��猇�ĿDh�W�]��h�0��m"�:�9m5E|�څ��E��!�e����«���=�����/8���z^��}*����{�Q�i�=[�3���"�_�d��|��</�q;�r~-p��e���q�!'M��w6�À��γ�l^۴E��z��*J�cK��Vݡ�!ad�@R/lœ̛\�q��zlj�-�p"�S^,�"���v7�L�\pe�p��t�:,3X���C�Y�oS�� ���?OVO۹.mZ��LG��@O���)U��z�ڑ܊�+N8����>yJ�#0����]5̙W� (<��Ȧ��,۱N��1P=��Z}"��!���x�9>����2W�قA�b<��	��i��@m�?�=8
�B7N�y&��eO�AN���Z�}] 4r��E!=�4�OU� �}�f��FW���b���S�̩�y�{#2fmtP���o^(e;�E�C9V�#ld���x96�K���kg��
�p�V��:�*H��:>���K�X��yt��·nk�`㣫���B�y���|���jd�k�ti[��N���A��X���>��E��"���K����$��e�����M#�R��l���"ۥ� ���^�c�洝i��b�<��N��t��u���5�ߍ-���A&�]i`=� G����F�V�`�ߑ�(�@�l�5e@�j��V%��v��Q��/�*٣Y���T�(�CM=��J�S�����FC4�poy�]B�����RoGDa�E��Q�Y�S��f��{J����ѻ�	{����m$����&V�,��w�{O����C��1�N�T���h�.܀�pI/����J�6 ���~�P�Y��|(����T�M&O?�6=�y�A(u��l�J�Z]{ Xn=ں�∪�� SÑ�7����7�y����V�H�Q7?�UZ��4�Ҝ���wo��<��X��1
����%�*xPW��.w�E�x3O�Z�	+��a���xg�0V/���	��eG��Z�RO�C%��d�V�,�g�ӎk9t�)�Maf���	��^�V��׺#���7��>�C�%���^��j;��Ɠ|0���^W��X�k[�Wz��T��%(���҂�9��dM�売��ȩJ���3K���$��h�;�X����d�v)0��ƼD��C�Y?lFv��ʳm��m���p,$�/͊����~TK�a��o�p6��5�ڶ 8��Ad�8���Y�^�.�����wwX���+Z� �k�����Q���y���b���+�5�7�**d-�o���\���	�0�]���>���śpC�%[�s#k�GF��-��[���I*�����)���/���K&�m�r���9�T�����-�iO��S'��������a��@�>���*��2�N�3�,x9q׽5p���j	�s�����O�'EF����-x޵��Q|ݯ����Y��ha��i�����,�OM2ȏ��5�s��O)x�{��U�5���X0�15��]P��t&m�l:���%�Ƿw,/&۵�E�����0e[Mߊl�	�I���T�U�cN�s�X��
���A+u�$���#����꜠�vi1U��מ�(׻����ɕ�f#M@P4<� 3�S�;�� ���9�5���:���:��yH׮9Ft�����ё��Z�����_��^p%q����,ϰ�s}�3թ�ƽ�ɳ����*��S�����,�!c??B6�3;T�f��l�r��}+E~B@1�	>i�7i�m�jW���)�������:�7�K����r�Eτ�^d=�7Б���XLW�X7���p!�)��0k�W�3 ��-ɩA$��N��|�����>y�z#���"j3��+\�Ret��Wa懯�V��DzC�ߥF�S5JJ%���y)�,H��`���k�c��5� ����y�r�<����{�-Usd��.p����k��'@�4rmy�R�$������!�\��'�/�MS�)�
y ����m�OS�P���D�>)x��"�
oB!_��T[1��2`�7��)��+�-!�Sp^ͥ�4���V�G.���h/�����;R�m�0*ؐz&n�jJNX^�.�l>�@����@�w�[���;�w_''o%��Q�i'��JN�_h{��m�؟bl�21Z�ͨ�θX��qei�53|�[	ډ3��E���)D�f�zP�;ks!�nR�ek��Yr(���h��e�����˭"�5��G�\����Y@uŀ=<d���m���i���|y�u��e�w���%[�@@��4r=���u��qf*��d�:�
��*�M�S�䦁bw����2������[�Stl�tm�s&DXb�>��-�[)`�\sQG�DĘΆK������Y$e �ˠ��@9��)��Mm�~���c��O�	,�B���tma^�CF..��A�'�Z�	��_L�m'�v�A��CQo)Y>�9��@~4Ǜ*C�,��aEc @Sϝ��`�S��$�O�VF��$��1�h�Ϧʢ7U�q(~��cu�<(~:rplL�p��9���oNs����f��7Q!z�6��¿�۞��fe�:�9�l�����%�|Lw|�cU�!���,;��q0��=��ܫJ>W$���u.��4;�šZH"���p���7)-�&�#��P��b�m+6]�a��2\��s�Uv��6��i�l����N�\��
����3Y�:n8w
ii�{��{k�<J���n�JH7SN^�0�(��/AL,:/�R;��ż���v��WBrO�M��s�k-1� D��	,�:��?tLYD�x�v�����Dy����rZC���@V:��r���@>�Ǭ<O�o��m�i���d���1���-Z��(���5�\��NĘ3�8*�bf�fe{��Ov�3@�(�����,`;�����{;ɣ�i� ��+�9R�d�ܱ��W�8�@	V���)��.�s�B��2��Z8�GÕ-�V끰�U|�}#���ԛ����ʥF
TIR}�>.v�MF�f��`�h �`�+*��#�ٵ/C��H�"�'���ǔ�U"{5U�� ,I�}�T��U�4�ElhO��&�N�������{9�4�]����*>��6:�؍Bt(�3�U�4�����,�b� h��3_���{����M�	n�5n�g~V|t)�+%ێ��ӢF7��<�;1|bIHѠ�s�V�� ��)�g+Tg�ő �)0�+Y2MW��"��k���{)֧�i��<]��h��jv��%���[�k�נ}tz�7o�53�9��|3E�?�'Y̹'�l���x�W����oI�A~%�	Ó?���#<�|�����L�����q׿�Sk�g�xU�^.Z���1�߼�ѯ�4���q)gx���M�`����P2pZ�Z���NR�<�㬺����5[�'�����[#'�<WĨ��̲���t��T�0��c� zKg3��R{/�w����^pQ #����"Zi2��(���]���~|��>�H�`ႍb[m��[��lv�ѡ�o2�UϋNQK���U������W8}� >ZW;��={{��T��4e)!��;�4A������V��d�Ck?ί��u?~Li8��3z�� 73����Exg8�a�� ���nm��>��Ρ ��������hR� I.�;�������I���£�����`~����%�r���>���@����_ ����PKZ�EN>���-�K	�=l�����ٯ�>�U_�� ��O�?l\1Xy�+pEoMn�噐/�0���K��=Pl�M�6d������~�«!�Ĵ�,�с�7`�;w/�h�'�����j�>�Hg����8�Sճ鏰�v��v[��<���]��D���Bx9M�c�-��E�D2J�/��5N�N �`�n>���JfǓ(��d�� ��*x�j�K���&�������,}�K1�Q�Z�]�ttl�F�P~�*\
G��0�l�X*�33Y���]��h�C����-�ż��शp��/c�(-�ޖ����."��9z�?owP�&�l�:��ez�U)�u��p����5��u��U��"Y�NF���v�`4[ǀ�$���,��o��Q�� �8V�V��bj=i�s���O�gվ�yy�<}�bZ�npO���nxQ��G�	�&o��	Di���gzI1�3����y;2fb�HiƔ�{�m�yg*��:�;�_�E�l�&���x$��2�_�ό�9�7�mqzi����=��)%��I��k>�'+�Lv ��'Bh�>�74��֨�i�V[��)h��� � ̞��-ܓ�~����f5�L)�L��~|���'���b�Z�¿5����g����TzRb�c�J��U�ZA�g��!����z�rZj7��=m���1�3�u�0����b��í��}��h��Q��q��Sn��.xr�P}�sE=��G�%��-2��[�ɋ��
��&NÝ�L�A�A@��j�����!e~��Z�òAR�1�8~�m��t��$9�_`�A �l�t�eH1?#k݆x~�S*�P��-�o����|>"?��Д7��pb���"�0��Lu
�.�z�vh�ةC��I�#U���Q�r�~�+���~��yu�,�7��j� ~�����z/�إ�iscE�6���ȯN������ց����pV����rXO��o>?�jp����y��X��`X�S)Ul�P��<E�Җ4���� v-�x�N��޾�XQK7��Pk��σ��50O��Ϲ�Ȁ���aC�~%�o��
?�8o��J�,Q�'�kg�@:�K�
	�	qa�f��n� `���e�jx1�}O�ј�ڐ0+C��ضH�������M�j�m/]�B���Ċ&�i�Xsv�t�@�=Mڱ�
}������7�pU���X�r^����U�9��y��uޡ��&Y*�W0p�v>��c����!c�&G���-A����C?S��<,���=�(�P��)W�����S��Њ�1a�Cմ,�Pzw詶|��B��|�t�����zy����VrV��"��Z�B*��K�v�9�w��ா&r��<D
�V�it@�Z����7O�����Þmo��j��}�*i�~:n��q��I>�=�Y���V�ڹ�*5"cc�}�^- �7P�ǀ�~aA�>���'/�����L��c#c����dw����	�*�sP���vފc�ȹ_w�\��q����/�l��;�	���ۢ�7gx#���GJ�[k��=���o�L~FGe]Vۂ����Д�"mE0e���@� #�!�;e9�6�U�,�����]����q�i�2���:y·�(qPWX�U�ju��?rǳ[��!8$U�3]j�h�#렑@��yn����^2�U��#��#9�z���-y���F�zoY�}�;�VR]oN�D�u�Z�Q�Qk��{q����!$���3,��.��!�����|<g?꩝

t��E{�"�>�%�/_�ֿ�ǮvB�g0`K������Z�=�<`�Ku�ѢGY	�ߐ ���C8�$�����`Cw�,��z�#�wA�� �����o�5G��k[�G^��EN��qt&�M�ӜE��ge@�JBi�g �|�#s@Q1�$w���YA�VG�'�}��ҡa�7�#T�<��ث6�MDv����e��\��es`8�z6|]���m���	�1S�::W}\`Ύ�N�����"��}>;�;!ڂ��n�/���^:����*E�s��ǡ.�0D��$�f���[A��C�;�Έ��SlL/V���~�
�nY��7=�����X D "�_������M�R�/���5���Pt��0�pn1��5d��ϺJ,K��<��:^�O�4�RSN?�KZ*�Ϧ�z�L#<g��5OK�9!�Q��s!m�V�.}WO�}�bb*e���1�~`��J$r�qU]�L��mh��/+9��`����\����Xs�LN\��7�[�c>H�2ͱ��V4x�;m_�S7hA=w��L<F�dj�	+v��H�@�D7����nҐ�������~F��Qj�8��|���|%���(p1��@Œ^���q��J�P�M+o|�z���^��Jk�g���+w��� �썖S���UQl���؜�!��Gx^]:zU���������"���^���K���W:@Yyf�%�y�p벯GȆ���!�;Y��
��l4{�3�|�H��s��#���+�"���聱(�##��;ۓ��w�
>iM7�֓ڥ,+��} ^߰B�d�.˨�-c�Ve�#'�P� �ۛ1�KnD�'�l�g�}Ï�Jч8D��`��	�����z���R+�;I�^ ���:AX:�(i�є �l�I9�q�,�l2C\�-�v��m@�|�f��HFc���ΰ3��?ϭ�&,��YX��B9C�'�]��]%;3��vau��3��*p��NT�=�>�IK��ß_�~܆�n9���Z�ׯ�}e��2�p�Mh?�A`wP��P�E'
�@c�}y�a�[��fYq~�!XL��L'��'�#��Q2W��o���kjJE�5=�فC�P"3���/��a~V���$�}�x�Z��V
��kZ�Qҵ�׾�
�� ּ~�����4�)�6�}�-g}�f�Z�,�F��DK�C���$��u4>h�� '��a��C��8SN��} sGTY�ᖼ�G�g�ucR�1 �m>D� t�\g6�1f�<�R^�^Nɿ|�&0\���}�3vƆM<���������CA*!�D���?�Ic�ѷ�A��~]������9�I."u"�ZI�� <�s3b��7�m�u�p��j�]��R��$%fa��9�h<�8���M��<�IA�̲f��z�'�Ur��wm&��m���Z���a	�E��a �z:Ξ��J\ip���(��*�V�0��n�wcOJOt�A�/�Eb �l[���8X��b�*d�&b�h���?^	����N�V�v �C��z���B�.��� a�j��� )q���'\� �f4��l�W���&XE��+1�ʺ\M��l��&�!!�Q����P���U׍�^�}i�}�q�L�RN(ᑸC|.ʆV�Ko�A!�����6�y��m1``�y:�O2E	��*MОؙ"��)t2j���Y@q$]��?{��C9B��n�<= O�Z�~}Vݚ-��a���v��`Aj�U+�����0nW�����v�b������y膯.���X�.ɩ!1Ԫ��@ඎ�
���O�u�<&X����ٟ�R����G���,��p�]�8�e\���I��i���GϸQ��@�/v������}�G��d�j���U��k��ʧS�i��zN��(�,J�>��y9��w�ͮj?�G��}ԄtU�rN�����Ia��%\2����ףޡ��j��Ȕ�����z˷a�#�KТ�����v~h"	g���"MK��{
(�W��k^�.���zXڶ�CO>����l���q
(�>�:a*�v�HLp��T;T�4���jA
,�GF�|��^4���J�$�\��fE#<N�8n�J,���\��1asא��Jv=�����zȼ]# n�eUVJ�����z|q��=P��N|wd��|}��t�і�������M���VWL&���6I� ��<�vi�����"z���u+B���me�9F=y-�
p�2.�?�>�z����5�]��8=�����סC݉�ē�١W@���%��u�I;u��a�N���xI�1�,l.��VQ��c83XV��{Z���ΰq�pw��h*��RA����cQ�y�����
z~7��$yY��7i��ʕ4��
���@ʖ]6��Ŏѻ3���g�l��~)2�0�O1���;�m��{���Y׈k�i/��g�՟�6m��������()�w6�v`xSY��X�Ƙ��5H�J|��~*$��QP���ڪ���9��#�Έ3���|Nd��z���D� `b�u�_�<����A�4!�?����K)��j�O������?��cj=ldw1a��ˬSv��HA��<G��ĴޛY��ؒ��1yv1I�&x�ǔ(n����%������{�Ygx���D[���OϏf/�C-��yJ��p�KE�����p����s-]mr[qf�A��krˮ�{�k��~���D�;���9^x/�(He���>H�Z���B$��[1Ql`�5_��p�m�ݬ	g..��O��?R�'K���'�@�H���׈M�C����eeV���\�������k�.{찤���`T
�\o��3Szh��9r�1Y[gM�ǐ+2�J&~�]��|l*��F� ���Ģ#=Rm��b�O���.���T�7.�W������1�HV�-��K��l��pm\���p텟�#vF�e�W���KT����K��&�F롐�&l\�&0躳�3�rF�K��,�V�H�x�? (p�>��P�IS">:	�q�)`�E<�kZ��dH~a���`�T��b\�LǴ�����R�y"��-\p\���s�KBGX�gKh_+�
�2K����q��k�7h�9JųMqY�I���'�����)Ӝ��m�(q^X׉Sy8�W��S)�.������F3�n��o|��:�s4�FolKćh�F�_l��Ӯ���{a_Ő�^�5,�j��[����v.�;-�B�j���[i�ï�X
��@U�	�҃F��n�bs��/i�%��#,��?�پ;��6���YG�c`OJ�ME�k,
2�朤O���Y�����@�x0���x��<e���fR�_��抵�s&�u�↭��f�gOOK<�P�ͅ������z8r�d�a�8O���4E�=���p�;ű�wbq	[�C�AC��CrrUn��[��} FH����˄ɥ�5�?�m�T�ywZ�?Ԟ���h�J�KT��:zַ����0�M�V��a؃�ӥ�H�\�K϶<}�T��s#v���7I�d�R��Uti�l(��uΆ�0+I���ukG���q5�:p���Aյ�j&�AD$�C���$�Z62ǣ��btЖ�� J��bq�O�z"�\�;����e�go�!d�T6�fW����`�֌~��~��PF�	��:�N��������lTkE�ďӪ�F2���>[��No�}kLF�<j�O`C�\I�^�V�a�6ރ�:��~���*$�I×�E�SϠ()(�+����o�U�3
�0�_3�?�9	:��t��@0O|��ee隑,(��n�7ͮ����s��L0_�P���[&n�����f��s��Dz�Щ�J��TN��g}mw1��_�l�ⵌ�O<�)��5�*p�@�t��_��ou