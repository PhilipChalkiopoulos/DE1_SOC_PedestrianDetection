��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b����m̈́��=��\o5_�K�	"������^[m�K>���"L�(��x3"��|�O�`}M	���)���e��	Ɖ	�G��,l�0���LDEQ��@|v���U��^�5����{�@{��z�Em�R�3���8���"��Ֆ͠@� �1 .����k��^��ur���H/��]ҧ�rW�}N�M�2�V�YX�����(�I��#��pNU�V�l*�V3C1>`�k���ϬU�=�9T�H6�Zd��X��we�j�Jl2�*/��a�tML n��7�x޽�?�E���%~��H�B�R�j-�օx�3���¶�⺄ǐ*s����<W�����k�N�o�Xq�@!>��8�F�C@i��>�ZS��W%L�����=��K���|uOI�&Nt�,�*��[KJ+�F�� �U�B[�F�[�tL�l��r�Lb���0z7�^��U�����"7��;>"�d{(�Di��4�Ld��_�qr�̯�q����x[B��]�7>��I�K����Hv&�u�Nxd�2D�W�h�\>奯HZ���E/	��!��dJε����p����*���H@���G!d�"r}e�˫^��,`���ah����2�e<z�%sa+t�y	q-
���}�r��b	����mc��<���b�8H��F΍�9�Fq����ш��[�f��(�mR6�H�>r�R���#.9�Y�����\�q�FI/9��B�ZE��v�Z��#���M��ݶ�i�{a h�����k�v��cm�!p]��YH=�xT{w~���#g���Y���.�eU��Õ_�$I䡉{�S���T ���-��+_ҏ�4�;�s���>�vp.����k`b����o��$��Q�N!>S�@��J.L���6�:�JQpňCEy�a0[�5L�j�$r��s4� ��9qx@��;�L�ˆ�7���"-����}3'P��vRu��I@����Z�{���*��e�e�� �J�rl�Ο�Hܧ�ѧ�B�r�����Cl-ao��Q�߈��Y8v6�u8�}l�#!�\�������&���΂\�_���)	ݒ��C�7`�.��������Z����<t`nF|�-�qG�$+1�qe�!�����P��
_�"᎒2�{�3�q�7�j��C���vj�h�+Q��a�@FWx�8CDv��V'Q�i��;��b8�1��"���@!��#�OA��+���	�2�غr-�1��K���>7�SX	]�80i���Zؕ��7d�&O�Lk)�X62�M9{��3eu5Gق�:}�ޫ�-4/��~��#����t����+��ק�䲕�Tj����E ���ъu�8_�*��6�}�5VB{Hk�2�6����	�.�ڈ�I�N`�ǧ��Hv��U+yV%O���38ƶ#@�p}��� �z
�����JYnB����![��C�rk~W
�~0u#���w��?��קg�J�XɄ�B���c\Ӂ�(�b�D��/䋉�WS�ȁ9�BHOjPy�_��(*�xl��o�@�t���"�ZX%N��V�t�a�F�滛��M�H�b��@������5)����c@�4=�:+�26	��1����I�k�"!��x�:����B� W#���6�G҆���,�*v3��4�����b�G�8�������0��y%�5j����Ӽ��Pq;�V:Ϟ�-�W��S,c��h�S]�@o�1v`e����<Ļ�\'^�>P$dMd /��pĊ�8X��̮�~q��Mk���Q�f�,҅ʋA�:����Ꜣ��/l~ߊ+W��<3�O7����rY]o�����;����Z��B���W>���n���\c�Mp౅��r���\�x�U���bd�0t�1�񁇺B��� �v��ԯF���K���Lzc�B�f!�y�Vtj�_��~�>����V)�_Y �z�nR�ţ��3�7��s�k��j=���&��+t锉3�C���\,����`���Fc�B�*�3Jۭ�=p{�S;��Uн�WC�S����D��G	�8(�h���ψ�mVu??��8����j��z��on�m�L����� ��m�~`���b��,�!�H.�����R��<��ꢨ��8f,�HV���W]���b��f�)aV���;�6Q0WT�w֧�g'ȯ\
�X�O1�!�嬭��aJ>c����[���<��MU��aBbn�1�F�V$rCk�O��8�#�a&�bq�W^0v��K���M�16�X����=�����d��kD���̖�9�n��@�E��D�|�eM� �6��"'�9�;-b"8��X��n��b}�./l�{�ɧD$�T��k����&d�������.z]C��}H�0����%]�b�C$���۹�&�|��flo���M>��Q1A�ԩ��
O����Ɲ7�j��q�5?ky��S��'��n�暋g�������ʁ��l3� 7��;�6Bǉ{B�IFоk%������R`I*�ET��6~�^LN5KH2��1V�gQ��/�E�ꭨm(�z�ֳ�l|8K���6����:�,������y�'fR�v��G���hC�&+�&,��tYI��$�CL=j�U]�=!R+�`�T1�x�1��Ej�od���s]ܨ������9G����:��B�5����ejd�E���.�0L���$�n��(y�6d�>���MF�H�5Hᖀ��DZ��O�j_$jl^_�/�\Y8a��0�oNL�O(^R�����v��S�~�u~�	�4�����ʞ�?���	K�˯�A:��W܉R�ncby}�,�`�.�Nx�h�5�f�()=�_Q��5�z�1���(���kx����~�\�9	�Y�G��.y��#�HL��iF1�N��A*ە���{z���)�!�V��~��۠�K�ܻ��?}�*ā6�|��NBF1��`��=�!r������1�d�޼2�^ �^��W�,�x��YJ�w���{l`��qv�A܄_���`��}�\�tI�&��c�z��7QF_����q�[��ۤ�ϐ�gZ�͈ 쿲z���Un�̐&I����Oƪ�&[/��($����O]�C�S}�h���/q}(E�}�Xܕ"���E��kW�W�K�������%k�A�J��m=��5��n�fxn/hn���}f��$N�`�<�z�������?������z���d�Q�ܾꡏ82�gtX7�_��˓���Q��Ʃ��6������<�j���vn1f����:�k.3��x-��/YħuAl9{4�hG�䃸^�P�TmS���"�Ki9%:��*_��+C���!� ��=l�m���cv5���#��g�^��$<7�0�&�RO���Q�$�J6�|�./�`��xK s~<�f]K�q�>���.P�V#�xdJ��`W���W��77	x���,��0d<�I���PG����p�����j���rQiAX�����=����ݫ�E~ �Z�:(]K�w�Zy^�\1����p�#�N��K�6^�ٽm+�S��r��z
ϫUT[���x�mD΢��c�ٹ}ة�������E�0Ku	dv��������/������ ��/+��߯��G&G�z>��s� ��Ջ"��W�J��$Ю�n�sOjl��N
調��������Cp�""\/}x�@a3�����O�gl�>B\��le�⺴�K�D��f�M�_#�=H�t��%Z�q�.������$����V-M�IX`�Ͽ�C4�����Y��dV��^�U-;~�$&�k��p�ص��&��V4q���4��|m$	�Н(�O� %�� �.dD�TZ撙�N8t���a�I�����@�(['e�����n�C*������P_��<�B���M�95r];!��Ad�V��=��ʧy���	�$C+Nc{������wV�6_�P롪*��z+B�W\ZS���Y��톿c��0�W�2����0y��`kܰ�ÏgFk�3�p_�/�4�����`�����C�T�^ z;���]��H�I�)�����!?(�z.u�����zp�1��� W�%u�`�Z�4����PJ*>��&��+tV�y`�������-@1�ru&��W���f$�9x�0{E���D�L%����@"(��hO�s+Ǔб���fH�_(�ot�T*x8�������
*�Ŏc�� �e��J{;�-J�˞�_J��!��ZIԼ�SOVE�w��H�M�<���9m��J�6�\u����zX�9�E�A�ޕw���x����O>���{)<:�OnԑH�p���
Z/v��m���V4۾ɴ%�x��ы���0���,@׺��Ud����Ơl���B�j������M�,F��:W�բ㘖a`I��@2���R}�_X'�,w��J�WyW�[TC䘺����]��dRTc�����![����������Cu�:�k��)�֜�Fd���9x�:}�u]�ms-VI'�=����1W����p6���[���L�2e���SaL�۸cӾ�~a*��ئ20c���M�-��/�&���|�>�kB�֣�%ξ�D�ja&Oq�&�����2`�e�?��������΍���>�_�{������D?V��ڮ'�:��X�@M��2���D��󴡅�,����I�^�پ+��l~�����|�#e26�&L�l�f G�ڶ^�z��~(��.r`K��2+�B�L���)MV�k�H���lj�a.��3Jij����E.[.s��3�Q�s��+D��2�ɏ�+&a���f&|"��+�Ҏt�Eb����r��;آ�0�q�r�jGR�Pad'���v{�d����'!��Ω��т���A���:�q�Cߜ��,#ozҌ�߂�?uS�����g���M�&��v�t���i��n��u�o^�s�-rJ�����P1֊���P�ڇ荴����U�62�M�V>�����=� 93�����O�DFk��/�|����ηfb���ʿ�#�x C��d��b��PT�F��RKV��'ک���i���3���( y�Y���3u��+�'*�e�`�ck��p$ ���b��F�8��\���� ��B+r���v*9�D���X���'h�!jJ*���svP�!<ل��"m�A�=h�FQ˷`��wX�ijA�H?�Y�k�������{��M��k���\]�=P_���*'� tM�ф@z/L6�g������T|��m���C�O��ԌW�eĂ��Yw���ư�z�f�h#���6~{��JK���N��7�`)�������:jT����n�lX��S�ov��L��J����v-{��6-��8�K��J �N��D+�|��U�!��"���x4�a_e�i��B6f�<�Hŧu���I�]�$��*��*�̇|,��	��F^|��ĳl��ǜb�ń��T�����L��1��'g��Cտ�=bnN8;�`�Ŗ����JS�Ӊ�ni��n12u��I����� `&���Jt��Y(/U ����� ��j���\"����-�XI@p#�y@��G���ޏS�,�f����4�{� lg��@�."B�z�~�����b�H�\�mHf�}�AjyaCB�aA\S'E�|���`�8(�}�.��������#o�&���kO��?J���j���<Y=E��n{8~ݪ�%@Mh���k��;'�5q�Q��$�������oT0�"�.�����c�w��Y�&�0�ʧ��. ; �����#� 1���|��F��ɫ�ہ�;}MYV6$:��32�]���(����A�B+5\>����k�g$[� tb6�xr1����UW9<�:��!8X�}Q��2��]�{�����J���g1/�$�d�o8��`���əKg�bǡV��/�	sG��<�fկ��z��4ϕ���q�͎+��� � ��ˁY�,��~,��@iއ�||�g�0cX��O��%/��C|����QA��%��9�÷8����[0�R^	J�EQ���fE�mf ����]����^�a�,P�lF�H���.Ǵ��d���ѝ-UJ~`32��>ͦ������w�zbGj����d^���<�4�P�ۯb/��"U����w��eT��ۄ��*�U�K:���a��~�Z�}�}�8	�O�P2�F�>t�+�k4��F��0=�b��Ĉ�(��h��S�������H%[	~��j��ik�,���(��[:([+�Od����72��ܳ���;{m��X��mE�� ����ak���8�+"biϨn�h2��J�A��"�c�=F�q�E�b��X}�~OۺAw�|L�[ꔐ�}��j�5 7f;EvU��p�+n��~mo붖D�X7	�}(��#���ѫJ�f�e��N`i_0Rҿa�����9#^`+��?D5�Z�t����/���pZ��r����}h&�����)L������/@�.��lo �B���}Wk�������+�QGV�L�n>@��C\����Q���2[5���E�?<��Hz�2�Pܮ���L�'���,]m�(�οÝ���$�cR�|���IZ�[��Z�s��|���hCa{i���p�����u�C��Jf�)�3{�0%v�K��]�D�j��K켦p�"� ���%�{�B73�uG�_�XL��O�F.Z[#�q��8��?�\��p�	���p$_���L��ҍ�L�����}���������.�r�&)����'���1�s�ڛ<ќ�p��\���V
�g^��CҤ��V��)2(~m�g�����"2�]a��� 5]��`.��A_��p����$g�ӵ!�ȨI܉FI"+��q�B��
7eI�l��@������$�^	�z<��+��ׇ��K[�n��"��81�֯�b�����}#g�~YY��rK���m�k��٭ќ�La��!��G�Č����D���o�&��&b�fW(�N�~*�_���ӢOܳf-Ф4c�\6(�
��9:7��U�b�ʜ��g�~𲯈|����������⠪�쀸�O�ރ���X��~o�'e�ZI]�E�>�M�uU_殏�T�Ѳ����<��2N�O0f��!a~�Եp*��YZ9]=�Q�J �����k�BGݣ��:��DAz/ͻ�.������0�tC0�����B°�w(0��E�U�J��9�\!W�?�v�9T��|�tx/>,<FR����z
E�,=�94�0U�}	�!&���_�(��w#SM"Xd�0��AT����J�V8Q��IF]�IVv���Y3>_#Hk��<-���s���ۛ?��L��*�r�����S�����=�>Y��tQL��ǲ����G�I3��?����A�b�RW��f'�-%�:��iA�nj���=�2A��]g�E��=:}�1`��������姱W�c|e�! 4Ӹ[F	�� ��=��+�.y,��]����Bg4�[���~~I��~���q����+q��!rY��$������kJ�-8�y�d�6�F�`�������2�B�M���P��ڎ&4���VӅ�9�y}���r����t��9�O��/��f�\���4�Qx1��t�aA��´�̯�cW�>)�t�M�í�Ҳo��Ü�T�6���Τ*�\����V�O{�:�Z	7�+?�I�,�&(J���ﺓ��v
��-ϡ<�Lӽ�왨�<�i�I��Gp�A��<i6'd����1��üUQN�ヘh��ɕ%5-��Ɖ6z��ǙBO�o�%�e#�p��6�|�����{W9^l^)!�{hȉ���E[F�x��vbxk��Y�V�� ;��~��5J<�pf�M]�D0����aW����!4~�d�Մ��W�8ӟ�3Y�uF��N{"_npJɃ-����y�Xoӝ|W#0L�\�`kk'2��tP'h��$r��f�L�s`k�ځ�Rn)t���L�����=�􍎩B�;�wQ�yq:c�	�P?��b��K��8Ϧ��Qbj��d�cu�RJ���٦;���Ss9��dςGP����)ӌ�x�O4S����wJ�s��`��}&(a=����$[�Qm޸2RH�K�R6=S�(��z����^xC��*bh;�+��3&��,x_�}�e�{�$b��ͦ]�A�W�W��Ж�:�Dr�7@����v$w����>z?P���o���N\�w�>3� �+��S�qLB���ꋊ�D�P7�� ��ρh.8�$]	���Ş��%�,���d[��R���F$O�w~&_X��)�y2� o@(B[�7�/���a��o��<���s�<(z:�Cl�^�~��N3d�;Ǵ!��X��G��Z�jt!Pt�0G&��}{=�6't�.<�!��y���k=J*�N?��~P�����;�r����ki�JO��/�&ľ��;�}W��4�}}%@�-b�-�O`rF�f�.�E�����?/�^.iꗥƭ���ۃ
	Xt1�n �PQ�!x`d�+�.k�UX}�F����!���ҵW���eM#s��0�w?�bA����su�@��j�F-~�a,�����c�dd��E�O���<e���g�q=<�O���0Qy���1��D"� 򶶵���w�b�ʞb��Y�a�F��y����F�������޽�W¡���kfp��ib���i3y��r�� �uo��7�x^�#������ ښc���tQ�6��Out�c,�h��rZE��m���qq����A?�E �?O�֧�=�q��29�2�$FL��x��$�o]`՟Y0�,+4�h����Lbc�+X}&<k���v�C�#Ԧ&kEM��˩����j�*Y�>,M'*����:�&D<s�Yj.��c��}��6���3g�Y2c��]�S��W��QhKEz3=�F4�V����k���wX��0��U�3"U��x�4��c�DpŅp���.m�d�������ji�
z+������TD;Ut���T�K��<�o��=H)Q�]�Y(�ug�7�kOJ#��ѓqЍ	�#��$�5g������Ta5r+�	G�QMɂc��P���n��L��i�SeM�u\Yq�[GR;E��V n"roR&t\� o2�
���sSnN+<��Q]�m���X���{)��e�7��r��?����d���k�+��*��3ޙ*���y胴Æ>�
���C�Ԝ_��%�����(�噒�����Y� _ZYicWO�`�~�(�A��Ҳ`��a� ͛|�Z���V,��8 ��q���o)�ٮ~/����(�f�ᙲs4�AnELK�[�).ڿY���=^h�5+�\���ǉC/S{������7���hb����v�
V���l��k[�u>�eT�Ȗkf噇��;_�O�d[��3�gnC�=�%1��S#5�zc�,x:N=,���<�U/�M���2^�ӝ<��-N��������?XF�L�N^�9(�^k4�0�_>���)�)}��<��1ګR���[��n;D����wpVݧ=����{&�<��[9�Q���3<���ܛxh�/���|eFG51��z>���e��5�!E>Au,��3�W̨׈�!�/��S�4\�4ki7�-�Z�H�Pa����+�v��3���c��Mut�"��kEF.~��|�
f����Q�֘*��˫,�x-`6�h�Ǚ�Q�\��+����
nmV?c��7 �	0^A�+�'����+�O_���Y%z�Z`�v��-L�����eyb�ئ.�9���u���u�h*��ΤG�(ʑ��p�@D_����P�]i|�Եb�ċi������6^z�����S�x���)�Γ%�?}xKo
hʙ�2M�6��@����E�˖��ñ����bF���>��k�:�=��_��9J`��?�Fl}j��ec���Axe��RX�Fܤq9���;h�0ӭ�3�4�eWo�j-9���[yA�(��[V��#^f�\��ŔӔ+�5�0�Q��:^�
�A[ ��4kGa2�(�ňz����75���L��_C���{BH3Ηi=��)<oR�ㅋ���ğ��J�]��f��&�[9�$��c��>e�7DO���+6,�L�%�GE�g��h�t�e�ws�&#:����g�Kad��ʄ`�M�R�3t�I�S���*�l��3�U�=�?���/LJ!vFڨ���7�� #JX��O�Nq�unDY({Ĭ��8څE�[DU�����\2
-+��ϰB �6�K�x�
15^㳉`�����������Th�u��&z��~�MlsV$�KZ����k�5��W�c���C>����xa�~#��A�g�w錫��c��J&_�	H�Y��w\���G#'���4&�t�����t���՜R�{׋)Z�y��5/~Z�V_�̎�,7%-��lJ8�p���j���;�p���r����\���b�pjF��sC��b7�5�����M�Utd�?P��)0��^~=�x5j������be~|�ݔo܃�ϙ���"��H:��
�>�@s�Υ�*�Dk�˔�u�ya�A�G�6��.*�r#u��W�/�k���"Hƙ�Uw��Hʌ#�4+��z]�.��= ���-�PU�g�Y�bq
|�r���=C��jj>�C�7�&%��>���[M9����������=�G���,�R~��d}��_i��fηX0�ҤG���6�4�83���F���3�����S�ӭ�Q����3@ʝ1�G�-�4��YO���������b���]|���[��q?������I�ט2�U;!�t������!�Q��z`;��B[q���ň�� iE|�k�k�Z��$iJc�r�(3�|]P���tcE��M �����
�v�࿧��@�mL%x���n)�z��456v���I�;��ޙ��*zd���D�͝���' �_=h��:�<6����PrX�D�����e�$�A�~"}�|�y��Q�5^��N�Ԓ�p�2X�����]�L�˄�]ϒNU���&(�ɽi9Yq�(����葞08��u�	��b�$=�Eջ�l�����`?�ˣ�Uf�^`�:%��7�(�#�?�Y*�_*�􂉖�k��.Z@r�������8���8:3~	�L)�l��|��a��J3�ʽ,v61�_FONV8x*��9~�)�<5RCM;^�hl�����ǽn�}��lwdJ�0�QP�sGKY]�����25�T)�PNU�z����=6l�i,9��9�����yPƇ��r�����D� a��ݸU���;$s�!����t;�~X��v}�