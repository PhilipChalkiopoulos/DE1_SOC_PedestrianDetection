��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z��4֬��9�A��;Un��Gh[�����<�#�L�-8�o����X0v�c�4��S�`U��� ik�{=�g]�C�+a
>kN}%]q�]���g��k���Y1��Ǟ�H� �a�C��O�m��݆��Ɋ�h݀Į��C���'�(���ɉ:�l}����K�fMm�p�����P_��#Y�aE6cP*���=`�̔�G�y���0��#��h߮�_�}�tW���G�êY��_��ږ:a[�r�KĿ�]^�[2_1��E�@�n�e��������G�(^@3�"|#,7��~M�U��(�����S��Q��K���X���s��, HE����7��I���'��?u���-�(�as���[��VQ�ZC'�n̭F�V��Y��<M��T���eN��$Q�Y�.�b#�|P�^�0�Ov���~���ߴ�A��!"��V�Ί��9�c���_%{;'Л�OE�e����~ɩ���~`�Т__&����"�J�R���u�+FV6����b��1�o2���BG-n²}g�C�S�	��ZZ�9�G�;\���C��Ơrܑ��$b��� ����;>m�i�~��ؤ��pZ�pI�_��u�[�B�\�Ӛ�/Ȳ��J���׮T��
Y�:LuND�CV�>6e5jho&{�א�^�PP���b�J��yP��@��v���:��A����D]�g���H�a��~*X(��щ�U���>?�˽����e�a (��J�ҶA�?G�_���PĻ��^�s�kU��s5SG҇S#��%�f�Мd�nӅD (�VԎ��_��(d�� �QF ��	�p�����C�C�L`GT�cw©i�Zh���)�#uI����b��c�A�{E,�F�O����W�C�KW$�\t���,�)�\��JqC.���P� 3��g7�i*vR't��ܞוӄR��Xy�7O��)
�/��,��Dr-�p"�]a p��eK�E�v2l/C!� ��I�ն��A�rA�+�C��s�۸,I5��q�����{wk���:�%�c�t�G'�|y�#���-k��p���j$��|���}H8��U���x�:l��1E����A&��vgb�:O&(=�Ʉ��\w��R͈� ���o\�@}�q�Fs���?j���rI.�3�C��*nYC�~�
l���ͤ���n��d������%bI$wł ^�p��0�`�/%𯰒*�Ǎ��"
���f�������|�=�J��5+Lˋ���������q$~�@�L��Ȳ��ĝz��uCR]�=[)h���VK�m����$���
(E�퀥2]�a"亦ϐ��HY2馫$��M�$�L�݊����*�j�!�o��|�WG۲�C27�ۊ���s����z��Y�.T�X�u0��P{�^���?^.��ۉ^�	�8\�a�ٔ//�P�;�\m 42c�����4�\Ȫ�dԧ��X�;oG���8����)��E	d����e\(��������P�y�`"��eXa˒�oݥ�3�J��_X�g�6j��$�>�	@��h+��������s��Բ��@��/h�Fʻ��J�%�`&ޡ�����sFA��J�C��<�Q���E�ԕuQ����5v�K��.C�
�����d���)qz���2�o?Y�ʗXH�񒘰3#"ya�g�Wn���jۥ6{k�U���oQ;*!<��ft�r�SQQ��rl����R����`��ڼd�9Bd�o��i�P��,�YѴ4RT��Φ�S3X��������_U��c��~a'У�GU?�����c�ݥn|Kn1�Z�wˮ"!������.z�w2,]�1�&ڍ;���S	�����!bi1�!�i�C������Ű�A��_��,���բQb�l�g;8�u�Xr/����Q��oٱ�|�.x; ���X�� ��3�o*XJ�N�yZ9�8��n�NPN��'�\�,Y�'���8�A6GxG`K=HX�y^��m���4��m���Eт�29W���J�3�����W��^dTd��7��@P��ɻ�_'�h#�ۍ>�>X��U�1�f*��l�~�Vz����+���r
W�$�0!G4�>���~���6l�c1��9GH͹�X�4߰���5�_F,.�ӠHJ� 
�n^?��T��@_��,*�U(AU�!1N�Q��,�6ے+�$Q��������H9P��|�M��b۩��3�՝���/�Ҁ5��)�UXϿ��y
�G�����[9�	?(�J�x�?ſ�5����?��PoD�aRr��d6��>��k*�F0@�X��f���sZ*��;-�9�[����S�$xA�9t��Jzw�(�ϝUVƁ9F��jI5�x��(5W15��z2�E���O6��M�{1����0���1Mx������j�c���'� �^b�9��F�&���E�NL�����tc�R��t^����1�s^��|l�/)�j	'��Al@J:���:�W���D!bSŪ��^͊�w�i"A�Z���&bGD�ʫ
�a5DL������<r����T��K�;ѿ���hx�b_����T�i2��7P�{�(κ?�b�����΢��1�1���6��6� ��%Wt����Cs�G]�9.�\9۳?�Wt�D%��o+�	�c���F�%�ReaV��r� �M"���Sֳ��j����3B���fIިp�5�c���W
�ˮ�
x{��_*��TC�d!�U����5�D�)�&`�����/[[ډ{���u�+z�#�ƶM�*wUڀdL�B ���4�; A�vu������p���)�:���^��ox���o�H���^��R�Iv%�{t�2��/;�C���|���|s��bvf|���踤��Iݝ�_�s�9�^(n!��^m���U��5���v\s;���J~g�1��*� \3�`��U����V��%Y�v�_t��Bҗ�P���5�~����y&2tS���տo����\�%�޳��4��Ga=|��9[������$Ө$������:���%��|++�p��M"?"�vV�a�U����{�<���֟��/Tip�9v�R�n:{G��Ci��Ǳ��4)��Qo]�2$K�h����$�挵g�Mit����0��EK����(y�+CF찹	��ituُ�����3.� j���8�����Z�����?���J��l�r�����jn+�Ŗ1'ӽn�Ü�w��M�Z������2샺��y>hd易����-��7��e-���A|�1�2�aK~���U�2�k��g�vxB	�Fh]�WNk�+33��^Ďa����@+�H�ȁ���{�
-r��쵗��y���A�tF�UP�
-�"ͼV�}��՘|ҩQ7	����������e���RE�<���EJs�(�{��.OD-��83�z�����t��^{�C28��c�`8m�[F�����ֹ�#�sN2���` "Ő�Q�;\Ȃ�\��Y�/� ����L�������aS�4�:�.ܝ��V�g�MƲ6������&��8!��i0(�"$�1+����ݳ��3�,��^�s=��D�i�^'���E�ӱ�"0]q�� ��IweC{iю�o�_���y,��D���,�{��-��� -w�/
F��> :�q";��F	�T�u+���{շ��*�w���{��}ˍf�O�\0�ep��=�V�)�����@t�%���)�
2�����|�9	+7�H=�sW����,�1YRD����DM���Y��M�����&�P���H����9Zv���r�aӳ�KY�g1�5�f��T�����m��(��Ú�t���@*�j����U�'TeD��h�.cM	m�X���Rޚ�(r�ܵ`}l��Ċ ����I1��F[�g����g5�]��@�T����d���ikY:.���LJھ�',�Af�M5�Yj�d��y�DVi����ML�� &V�p����t�<�4
��^��)���`R����y���*�����DTq�� �!��Y9��k�K��R��p��d��
L#ipf�J��	"v��QzB���FZS���px���uW���-65����oG:��V,������>�i��Mͳ�^ N��w￲xt�'��dn�Ϊ��Z��߅�(��B���*�B#����X��J��D��JA�@���G�uuH �?S�=�m-kʘѝl��Dv�!5�R��r�eO����n��]��o���Y���{�E����T�,<ի/Fc�w]E�	�L��6����u`���C����o��+��6�Q��끸�L�i)����K���!:V�����r'e�pM4ϊdXF%��s�u'[�ּMk�������H�'�x�냳S��y�I�_E�߽�_\�dbIJ]J$XYLe.�i�b�/w�*,�	���*�`6|gmy�{���������C�ӶNp��!o�j
eh��٢U��Xۘ�<h�,9|�y����CWC� �E# ң�=��]��C,��R2�U �A��,�]I�x�d��F�����l�P����(��f��~���gȽ+��а"�����ڱlJ���8L���{���vCץ��u�Z�
�A��۹ܖ�n�<O�Dk�YMlɽ��{��~�^�U]WB�t� ��2���EE�ӆ�TWr<e��p�h|��jqjv��c�NsZ��1��G��"CRR��(�I,^��_����-����Њ�����D�����B�����g���x�c�`�1Ś}L��&�~��� �(z��{��g�d�)��B��I DT�D�u��`��<��eב@j̇W�!��U,�b��0;����L�߁�2�N��S�85�&��=CX�
mz����7�o9��i@�cs�yU�by�����x��u�����i�XQ�gyC�E��@?�ĸᬤ˔2<�3���e��u����]�X�Z���n��_f>�������z7]v�-{�{������l|.�"i>M�7�'n�܊�Kd5(�`�Ly �_If;��U{Ӣ��<���n+u�9�|�x�����g�dqSЃ�|�8�Wf�A�Z�=r-��Őy�P�L�k?��+�A��c�j�G�[����k���f�C�F� �ᣋ��	�l𷥂>g�K�������KV���'���^�@�YT?!����g4<���iƧ�(HזB`�@�mNs�v��_Z���s4!��t���\C����sȞ��:,�[VN�3���L�73:��ydq�C��E0�,(J��^;Oghu��ߏ��v*r�C�a{��~�P�R�Ifwx��97�6�>����n� �����{�v�M��(H����~ik�<'B��j�/��ǡ�=W��JU�E��0���]�:̔�1[�6��p�����p�{}!�!�"}P�0�|�q�����Z���t��\�V�p��af�pK(v��'C��uf����4&��`!�g�p�;r]�oب���o�}1�5��h�^���V�ʁJ-��N	W}O|�C:$����I��g���Es�%Bj%V�M�Z���ݜ&��AM����]���	����$�t��L+����SB�~G��#��@��9-�$���_%��3� ���i�C`���^���Z3G�4�G�Y&��{���M� C�4�;�V���ذ�3�8~=�>o@�{��HොRX+@�Uۊ)�/7��/��=sa;�9�RPw��d�G��YM���B>(�8vs�V�h��@Usm>���g����y'�q�ֹ凿؊S+ ��M�E*$�t�m@_���|����{��~���t�U�3����c��;Z�{r%&�8ɑ�J��OĔ�+���ܔ�n8� ��P`i�r�J�P�}�����m����ĭ��K
�a�p�=�(\DQ]Y��C��Qe���W�J{�0�;���/`���M�b��wA�;,� ���Xq���T���dw� 6�Z�-��[<��H0�'�iyA�)������;	 mb�U��e�K�}�p�#�E���"6��Q�\���:�|��]�|;�ea���B���1.�_��]i�>��|��qb�/���;A��E!ϵ�,�h�ᗶ۶[�V��v69w��Gud���4�C��({jR���j=3�k��W��@!x�߲�D �ɸp��Q�#͈�,Xu�����$�6
H��
=ܥ?��l��%{����N$}���ޣ��PP#l�9�W-��b�j�������J+�������A�g����e
��]�BZ4(�Y�K��V7�,��њ��'���[꾚�Y���l�|w�Xp�Q�ܮ�\XIEx\�-����\�wq��c A�%��
��.QmBޙ�P��E�U~cJ�F�m��a	����\��H?;8����D�3��:z�5�09��(�D�g����Gc||,���T I]w�����w̛���7��jX�8l.�ѥhʫ��Ȳb����(���וl1�7|ǼӨ�+.����`b20C���j;�3��F�=1��g�zN'�m��,��Nw�؄��y��)}�+bǙ��%IJN#�?�һ�n��r��O����]��>�=ρ���^�rg4,jΓYH��"��@��몊����V�K�2
T4����BWCc���R�>gI�#�����u���w�	�nnB�>/���W;��$�yCݚK=&���1y��L�{�s���.�<󛭖�L�k��������	+��g�	�۪��R5a�u���ePӓݵ�<C�@���g��΍7������kI�,��[�݇�!�(���O��ɦ�i(u��.�뤗�^�M1�k,�1 ]�M��=�M�����*���v_,,4���b �e�+�L�	G`��56𳐟�Jh� �:�� *O����兡.8��&�Z��9w��}ۢ�ʎ��}£pbP�+�z�����7(�i:��_#^#������c�y�ng�_pO�]Va�p�X[�E����g i�����R�U�i��?0�w���փ���}�� ���A��y�����ЛB��H�]N5�G\�]U��oC%z>�Ş_���r�H���Lv��O�`S�@.���ס��J$�窈$<-��\U�<���gD<�
3��]�x�ǡ!��"|oe(~j��-7���|�[0 �C��["���$�?}�b�s���p�%HHuYDO�:V��kݨ�`��&��Ɲ��yW�W�H��@�G��������j���q܃}:�8�r�����w�������O��Q7�椊@D�nɶ3N9e&�7��Z�.��Ӏ�F�7v{��D@?�B�C�O��=;k۶rKM�B��(C�,a\���8 ��b��=O�����F+R�%�ܳ�Y�ۅ���o���R`�#)�G�x��5e\pl+L""��L;?H��MyhKj/������n!�6�����psc�:.�Y�/���xٿ3���E�,g�^��	v@�|'W=��2�y�Ф�S�W�������[���/�\<��`�f���.z��<�1�R��Θ��,�:,?���|��ۏ�ϵ�1��<j�-E���Ea�`X����{s4��?,�`���CGS�Q��a�Di2����BM�q1�b�B� V��X�u����a�Ս�+}�}���������Z���7���:TI������ �G$ /��aT�*�R7�r54�n������Bd����c��F����K�����Y�������u!|���O�(�q<��t���@���Q����ge��q�2������-��d8��hE�؆L�޾n�!+���kҌ�|�$E��[�T'��֗����X�U�7G�2��h���#8��i�3��#On`ˤ�ڸ���r y(C�MZZ��+�����(�Q��)��E�TOYwx���/�f��/����M���t��l+�?�������Ӷ��;�+g��Հ��q�a��Mo������|��[Һ�1�������[�B�z�BQ�6ŀn���_#��|�	���Ŷ	�������}gxAG�A��'�[Z�%�ԇ>��X���`��cM�Or�)���c9F	�c����w���[*L�F�ö��^2Wň�7��S*��kӹU��Z	ԛ�Q;��̓�͢X��s0�,�:*O)�b���o��"��]E�m=8U� T����43�}�CPu�W�|��b9�X_��J�L�=wJ�m �i�e�C4P�G*�N<�r��?$ɻ��C��#�V:U1(��H|��ۭn۱�4n��G���]u2Ƕ%1��b_"b(��_�F#�P��0��:�u^}�s�N5����9��wm�ş��H���0��z7-"ʎ�oe�>u�`�{��e��B���:�}����w��WvY�j_f�#��k��M�n���x��tdb8Ue��+��/�h��e�����t�S�C���aO�� n��^@�I���rQ�hXD��ޜ������mi�[��p�u�nZ�j�Qm�iN����zV�'6�D���;��� N���U�1ק��}���'2���LU�=B<��Kd ���ͯl�j����=Ƒ�ǖd��^��N*˭��M��&���I�U�n�*�w�u�����#ɖh�=��H!�*�ܫbP��!�C"�.��╔\R*\�x`W�a����[F|`z �kH�����~��2��$y���V/	��_L��GT�Һh�_z�nI��nqբ�D�B�m!q�����w�g�ɞϨ#� �h�������2_p�N�Bk�̹ 7���8����Y�I�Lr���O�R����7CZ�m����ҥ3�����h5��5;���u),�i/�����6.)��J�S��f�}k m�(�/{gDJg�_�E�
d����S`O�&����	��
��O�g�G�i'!�ă���"���"���^Wei�DS��!w���$K��z�+��mY�.򱵅�;�V�vjbJi�Ï��D�Ʈ���"I���F����h=,ľ3#��(`�a��BQ�fBTL"��9��#����\$��\V$�&�4�&�X>��y������6^uWj߭&�[����J���Й_6�Zl�C>D[�@���2\ƒ%Ei��P�w���4�n|-iA�W�W���+o��v�7�&��z�+�X#��8�芏Ϸ�&��u=T#�_�K�/΄�)�f��ø>��N�[
_���G�#�S��I,*�=��H��U㼵���b;rI^�>�&�>�hfdǿ݅��ř#͑J_�?0��c�h�M.$�T��l����?����}��X)��eOz���+���f��U�0��nN��	�8^?tsPҪ���Z���5���G5������q�ކ��_$��ɿ�g�s͉���s`�f�ف�����(fH�G	ж	G�y�Q���Q
�~�0�|߿��H�A��e0YS���j:h����Ƽq2���$
���ߓ8K�<��}f*���	�J���^�xY��	&�5R�DE��8��_�{�o0/L��,��gpJ�;j(�e�+sHw��������;d��*�[�{��X���L���8�]b��WZ?�t�;i��vxl��t������$��>�����aɍkW�,j�=�E���8���_�Ÿ;���Մ')oS��bwʇ<(	�l�kP�k���Em��8i+���c	�c�S�r��a+�����v�U��Q�5��/�߬W�6kv����ُ$�7xo_ι��p�%��1�^�R`h7�1V�)Ĝ|��4�c܎*�v��ٽ�~�C��y���n������ ����~/���:S���Y��7�mA�Z?�f�T�����m���� �����*�_�!C��'�L�cs�u�iL�����T��oR�U�y���Ő1R�����;)	*`YI���m�a�nFF�e����*���u<�T��O[��
(+MJK0�H�=���4�K�{�"��{tPY�s	h��W>:_�V��;ͫd{)
=S7̼��
~��ZV�8<9�W��bv�4�a:"�S��u�s�|�=�^M�#�΄�R�$LW��WF�o 0���c��
�rf�6�ߞ=�ܰ��TJ��Z��F�k_�:v|�bn���t�����햼vKs�K��y.'cK��/���%��Ǥ�?!���*���(K���D4�!�B��
en�Ԝc��O}3�Ń(�v����0����6Һ��]Z.�1�c��4���R�g�r�Ͱ�-�v��h�;�ӓC��p��g�d���o�٭�I�V&�O���|3��༃�ON���As_�c<�6�r�m��n�8l�9�FG�ȧs��³��q�7�ۋǈ��^�� ޒ�q�#�������TtV)q�`O�O�ɇ���N�L���Yq���3`J!i;��߈��;x� ��f�c�~<�<��J��+����R�,�_���!R�=6��=^O����n��^�k��V���Uc�lX'�Ǆj���d$Z�'���֎ɽ�)x^��2�m	�����m=��@,9Q�M,6f�Xd)#��DEe���̈���-�맪6��Q/}��R"dE�*�4DF��[��OysU+UK�e7;׿#�P2�R���9�ҳ:�֣z�B��?M�tί�5l$�/��83��y'�R�Fx%@�<~��yp���`=��:=�+\~�X$�D9҂?� �5���i���(��Ȯ1��?QM�S+|@���	�oD!)�b�=t��"+Z��#����I_���K֨L(�����E�I�5�;�d 
G���q���(
�o5�:��3}$���a�S��� �>"�V�#��02\����m$�
L��f׫�pw/t�F��>%�m�#�#2�*��L���'���R�f|(�	�@	(8A��#��cp/�l���M>�#��Q��W^2yŒ9�IL�W[Vy?ؼ�낹a�c�S8f,��G[H����M#J4ÅC�[>'V+�43|����>E����Vo�)�V�&�Y�/�ap˔��>Udʤ`�\�wM�BUW�9I��iN*�Bś<JW�>����Cϑ�;�s²�ʮ���L���U��H�e�dW��;�]o9#?:HS�ƒ������u�#���0b��R��YB� �3���*� *���������&��\W���n�d��Q�3����Aa#�i�T|���w_���N��lւ6�pSR���T�qx�OUE��a��ɩ>�U#&�1M[&A��W���P擏�A��x��{%�Q|ת�k�3�r�+ �Bu*����y+y�V	�l��d��+e>Td�@|Ғ��y��}XH��7�:`���9���H��iX	$�9������_�NA�(�r���ye���H���.b Z8_�ĳ����ۍ*舺���,c,
��!�Q9-q����}J,V�!�xZ<i��f9�J�2��Drh ��"tΑ7�i�:�����%8�Y�ݔ��!�e�8�sE�����&Z,���X���8��oP��a9ycX��U�"��Wb��Ɍ�T�0�1JS��)�Dk�ߵCNCԷ�!=~�5L���ڪ�|O��PW��{��]`}g�[���K�LQZw�̿)�|2F�����d}�5�}�T%㐢�VČ:r"�*"arz�a)�''(�{��w���Ϣ1��7z&�מ:��\$\�ӯ��R�������@�A'��ܫ���Ehj����E�q�@2)����iq4��c�RG>k��h�0wc?�����}�[4��������Zg.%��ic�����<F�6��u�Q{���
�V8�DÊ2��3v���ɢ�eH�*�K&��0!t���X7%.���n�g��15�=��Pl'�+�<�v$Vrη[�?�񞥢�M�&	��y!<�hy@?4�?�#�rJL����|VC��(�h,��^I���J����p����o�X�x��ܛ���"[��茊��>%H�6��j�
��Y��c|y�2j��,�a�T����IsH ^���cX��S>�M�"��Z8�j	+���89��G'U�N��i���1��H�������f���J��������q���K9|~?��W ����4��� �J�J|�X��P�����=�K������x�{�����uMu�Y^
ܿ����x;�N���M�OѪ�-gLKzէ�~�wW�G�"=E����8H��5�p�������J���c��ځH�� f��х�,�[o�"x�i��+�@�=u�'a��o�(� ��sLn��Hq�U�c����S�g_^ʙ�Y9��-r�B�o)����;��`e�x'b���	ܠK��kr��~.�R�J0�^��O^��4�Nr��?��ܚ1�WUȋ����x�#cR�?	�X���\&7���Lt���ǝ�`O�2���{9�(_h�;�A�g}L�@d�y>�(h��~�]9�����Y��=�+p�CF��'�T��`��]��rT���~ ���O;Ĩ+���^hؗC�ė�,�r�9X��&�Y1D}H9 %���*�ݬy�@�v`GG��V�]��gU,5r��\U|��Հ�=��`��3z�t�e��~�	���d��J�	[��*�������jUj�,���2��zTF����)��%�7�-��d��ܖ�VN���|7���/d�0�d���ٮ�g�+����.��?=�>��vA�	�pG{^��(�-H�̯Y��l��h��Q�)܉������p#��<���Zt2zt��+VW};ٿ������Y�s$4U-�����w/��Yl%D0�H�ǿ,�j��]�R�W�r�Rp�1�*)��C�o1jm��Θ����%5�4ED�gxm���,��~@����?�k�/6L�}D�K�����3�O��;\O�6�9�#��V���1�O��MW�í�%�lK�%�	��������T�:�ѠYJ���тgL�ak�)8;��mwk��TaE}i$'&��u��,�+a��ڪ�%NV�E}�������Ih�#
�¿�',X'm�H���Ձ,q�TQ��������Z�ɤ�2ߜ$5�8HZҟH�Jp0���Fk���&`���0��M|���|����ƀ%�,�8�?��(��P4������Az�ybC/�=�Y�͏�0��%|�U�	�Cd:�[c��b�bȥ~���{[�ą�tr�H?��f�} �ݧ�e1�r�J%m��bcP�=�4�Ôp�aQ�~U�ԛ�\�vX��'v��,�ӓ�<Í�Z��l��E������B]����q;M���׻jO)�6ù!�����V�Jp�����+�0<���̽+���&��k��i�ߓGĽ( �idg��D�����(= "B��2��>E)+�q
���p�uS�ɔB��A�H]��z@��u����k?�w��� �x `��w����G��U--Z���f2�K��+��Zr��/�)#`>�;*�a8h��$- �!����t}~,�ٙ:�Q���:B|U��sɿV�K�x�����ی^| �YzL�u���?�� � S$t�~s�C<7��L�/K��W�?�ͭ8Z�T3��Y��<�ЍJDaI��Y,q�l�V�}c ��?z:;��Ϊbj�ٹ͞#$��F�D�rQ��
�4�`v�_b�X
0�< :׫h���lF�ni�7K��c���?����p6���j�B���k���i�"���s�|&ޟ�^���|���:�2� ����kt���5���G��Ө��NΣE�#�L��x����[��b(W7���4��~�t.x������O���+��b��r���F'[�]+��4�b��#ڿlDA1���Z���� ��2H�n4�O���w�E������ݸIj/k��TsV�C,R�KK2����v ~��߭��"K�6��Pa��o����^��|��F����@�j;�J���6|�.Tl����W$m���r$),��H��]��.��B���ʏ��QEi]�?���tt�1��r�]oޥ��1nD�3���v�sΥ�$q���h;Cg�/�
��Nb.���f��/]�O����#^��z�8��������Yg5�+{��yh����B���g �n�{Eb&���*+��v��5����Aʃ(�ݓ�� Am
����3H��7l�[�ot�x���z#IլR7����'x�9`�ڡ<,.mB��Z�o���q�"���qn�f�)��Y��r��wr�c�������+�9�)���\��c��еO�E�0�B�}�oq{��2�V��Zv�����qrP~6����	��4�`%�!�@�|W�Fʅ���	��9�8�����1��	Aۖ6�%�d�D��~�\�<��s���
�~��X^��N���W�؉v�u�m�7���%��*w(���҄˪�ZY'y5s��O��i��@�ԋ�((���$]bLS��)��j���sI��s���{HOw5ck�xI߄������� pT]Ny敗�AbD{j�[�&������Vؙ���ĞN�J= �������7Fa�83�E�����F��U��>��etFz��@����f8��PM3�:��3���s�����҉/���R����B�:n �
�J/���:����ٍ�5�X����
ǙHH�Z�D|l���^�r��iυ�Cf|��K,V�;D$��B;�U�[��i�0ms_Z�e:��\�X�*Q˺~92�s��-��eu��rN��ĥ��?(o�y�ݰ��I2�!�RÈ�����?Ԝ3/N=�!.���N]v�#�"�V4�b������nrPLcG�}L�o|(�Ń�ǂQsA�����.�a`�y��x��O���T�2�+ˏk�'�(:��0�w"˹P����
+؞;��E�h;��_ϥ�.×�N&��������Qo%��� w8���%UJ�"� G�^�>rƋN�b;�� ��?�C2��P�B(cGCwA�E�jN���Z&���	�G�D�4�>[��F����������� �Z;Þ1����B	���)���n|�/�����b�C�)���YN�N��%7C�����xTcfA4���[䥝w�]:���`by{,�{����lX�Ңh�Z�A����xa���RuS�+_�/ W[������Nݹ4��l���_��~ wIx6�層P�X���_� ���G'G��M��A5d�&��S1��_�(�E�l� J���ƅ�����SƯLFr N���5�l��(6�e7L� � #�G�Ġ��;E�C���[Cj��Kн����-W#�G:�����F�O��[��a��m����L"�<!�/��e�9+�	_����*Q3 g�O7]Yw8.��=��'��H(˞��q�v`����y)�����A��!��䅉UkU|s�fK��~�}>�t�E���H�C�r [Q�.�U��u*a|��/�)0�4/ƣΦ'��*�oo�H30�#t�Lu�)��=�+^�,���!��vW�q������>^�����e����~^�C."�Q��!�:p�yЛ��������G��1H!�����D�oC0�u�η���͎q��<Gg�(k�tٟ)0��e�U��km�K�#�:"�����8;�Em�tq�TZ��O�H�W��"oGtv���G�#z��M?���1o��^̪po�n2��'N{��Q��R�b�,�8��ja6�o�c6�q�x��J�$���D���Ya9c��Rv�����y2=�v�?���򯙛&����I"��i�3[t�U�����0N�υ��s{��Ov���l�|~�8�Ͷ���b�C}�w�e6�ۙ9��8w���n����Z(�PؔR)<�r),�ϊ$aU �[���]Ʊ��"x�{�;q��x�{�\��A$Tz�W,�;/�+�N��������Y:���Ҥ���ԙdG�K4�rNH�Ś��I�s�1"Ɨ��,�z ��#z����'�'����\��Z�m=����QZ�3.��������~��BDҊ�P�;w��$��_�� ����p5.,G{�ܞ	7��}���$L����~��ar��,��_r���F�L�v�� ��k����'D��k�?�'���R��C����L?$�.y[A�C���-�~��@��ޱS����?Q&���dE���d��3�/���h�V��b�����D�=��$e�?r&%��L���n�ޖ�đ�����6Ɖ�`Vǧ�c(�Uy�*K�z֞���T�S̸�
�y�?�?�_�%}�$-�]6.7���sY2#�'\S��p��ݿ�Xc
�u�����+��;#�! ����+�g�R�����b<�]���#.o`	`M�(���Oa u	u���Ǔ@�1���^�x5��1���8�w�g����pG���XmK8Mta?�;BD���o�`!�ØĚm&>�2�ØaJ,9.��9"�q#m��3��u����dO~,�k��T���x��Q���(ٺD�hH�������O���9ڡX�o~}L�e�����d>$�z��V�����Y[l-B�-�>8M�wG*��ŵa�'�n=�+���M[�z�n$uG�^9R�N	��$AC~.=�H�wj�s���Zꂂ��������u-�C���$��(<|I7 Y���O���V3{���k)%��%�^�Ɗ�T9��>�1& %���/��o�
]��BԤD��]�C?)K�{A�������."]�l��z�\k�0J������u�}�)�M��Ü*�_�5�����cXu�z���xL�̃�/\Ĕ�\\?�W�mcOE>��z3���2	��H�<O���D���[QE�̣p"h��%�_6L�l�m����$�[8��Ä���|�i���-�Q���9e�Ȍ3obɈ��Tpr��F���
�ka)�O�:�sT�܏��"��Q=+O�& ��]Ԝ|��]����A��]Հ�t]6��-בֿ��qvT��~u�,��L6
%a�L:�[��e$�/���#)��9�\���SLT��TD�,cڣQ��c[�J�a<\�b$m�);ґ��9۰�*����4Ԥ���Z��*h^뺸��z�"�:F7�l��g���/'�w�i��r�;�[�T�9��|j�wX�q$
���0�ŭ���V5��g:�w�����3�""� l�Vh~g�+���u�.��{d���-���q�_I`�l �Y�l̈���]���?j�?0��w'f~��,�M.��k��iݨ|���l -�Y����_ߒ����LX9�q��b[g��&��H�� ol
p%	P��`8Ir�*��t�n!~X1<�X��g��7V�O�{�Qܻ��S7��Z��U�b)�/�٭�����*,S!0(�y����6��^pK�(�A�+T���w�\ܢz[K����MŹTJ��v�4�=K2[@��J����a�r.<�A!���䷞���Jg�-e{��WE�"��Mع�'����'E���%ﯥ67[�*ְ���"WC,(�Y��~"!y�*��r5Y �-�����y�s�Rzo^B�QDͨw��$�wB}ǶU{��|`�3�(m�E35��&���=൨� �S'��2�ף���;�m[��ӧb��@�;�r��c��rPQy\�g�¤�"iR��"`E�_�~+��N�T�I��(v����<�i֧TN6�������I12�Sl?���M���t� ���Y���P��'���f��b%��H�����vd-�{�8�P�qQ�O![�l��c�������J�/e�s�s�K~8�������":��Lꛀ��C�*�~n~�ʤPN� ��+�������b�m:������}��^	fA���ő�&��=��{��g�<]� �
^�|$��=�{5Mzw�U�sTK�Ga�����F}�>�PSg���k�'�t�e�@u���2N w8ns��~aрQ:�CZ��j�H��5�������U�Ȩ1�e���&�Q����r����obh��`M�Klur�N� �'l��[�'8�*��?C�Lf���S���5/w��ϲ��K�߈�>������@�wǶ`�6������� b��uEQ<���y��p8�B������m��w�y���k�ו��lg�Q�4����B&��+Z���o����%�N����I�$8��¶��ª�2W_<n4_`*����xƢ$b~|$�p�%"�0�	�V,���"���F���+�	I��#0�y�|xKp��޻:f�r3��&��-ɀ�S� ��U��Ґ8���y�����|$�~!e��k*�_�h�u����%s�i�{0�ܝ,�ж��D�2�0�zS���G	��T�m��,E퓧������W�������� I�R��H�	ٯ�5��ں��4�D�;�s��+0/4�ܹ�pV�u��mK"X�Ys��i���K���i��Q��zKL{^B�ٸ���%胵�O���C�'��)��i�^A������ �tq��埪��9�JC�⨔8��N�J(�z��Ub�����g�MZ�_�Ŕ���|М�̓��g�=T��,�P�QI�/�É��kA�+��d |�����[��?�-X�s)��aW:K��-�Ǖ ?k$��h�&�|&�Z�͎��3vYE��7mz���J?��d��V����z�UX<x��:�tkb�4��"d�-A�m�V��'=v�����{1�|U��yi�U[O�"ܘ�{�N����x��p��ؙ�u^G�"Y�qXWWLd�dm4��C�z����?��a�ɗ̄M:š\��0����~]U��̀oG�<�_�.Q�:��Zr�6%�;N��]b=��N͈\�E�@_VJ݅g����PR�=A� C�-ɳ�����䊖����ʰ�N����VG��m6�c���_����	SZr�H�f�Qcu~@f�ɰ1S{L����e��@B�}H<�Ɍ}��}Y,���B�m����lz��an����y&��^f��Ӑe��BxQ0J��_p�osұ5�>�߁��ϛ;v���r
��V�QQ���-���Щ�#\:%�os���x��i��i�!zϡ�/��SGf�Q�в�x�������6rR
��.E+�9��y)
�;'J�O,|�uױר9	ꗂx\��#��b����D@�|�����粑9��M7��h|\��ù���5��O{��W�|�M?�~�L}��<K=~�[Hf�x"��!\��IS9��r�*��1�w�]~��w�sR�=��AC�W�hr��H�k�?��1���\��\\^g]}N����	�+O�eܽ��pVܪ�~��g����>��ؘ	22���W��H�s�|<�gU�;hK/��Q���ķ������Sb�.a(IW�K�Tw��`�Ƙl#C$�\�����<j3:�d�2��߬{����
j!��Yud����+���(U�ՒW(���;o����"�8#7�p7Ҧ>��Ҫ�������Np����#R�)�E�Ȣ��e��7����W��ks��;��2:��)�ɉBsrw��S��_�ӹw����y>L�/���2V���4�^�<^�zb)-��|�-"�Ҝx�fL��z�/ ��#��<�@vV	�2��B�ʝ���^0T�����'���oՄ�l��<��uޒ/P����L�T�N̜��֤��:<71�)�1�1���]���KCk�.jq8�F�q�n��C��z��rk�l,َCSDUB���{&z�{�6w�֯�6/��c�^{j>.�ථ�>s;�����RR�*�@�1oIZER�im��W4��2�Ndvv����@o�ؚ�D�@?���c���.xr��.h#Q5[�O	�M] k�O]0�VxZ^^Z�n�<mV'$~����a�'B�A=���R�"C[3M��5�Rxv�j�;kCu�	8Id�F�%�~2��&�}L7'�-oG�]Sͦ؍q�L3�o�^�B��������FAm�kp����@c�3hS'PZ�����~]*E5��^��5V �8�i<������~h�K|� 	�� ؆=ϒ�y�Q�N����򅷊�Z1�G��;���L.��g#����J��n���M�	����t~v$�8��]����>��֬D�Y�f�I�h�Q��@�bN�cW<��R�������iD1�`ه3�Rz�sG��x�W��Zu軓�����X�l[��R�����[w������2-�����Q�@��j���W1�F��;���Ժ����g��ڰ	��RL̋ˢ�32/�C H�Z�k�Fs0(=�ݶi�����0S�yvD��� ���'�L5"���e�+e���<{t<e�ᢌ�[�6Q���m��Leq��s�����g&F�~�G~��#���Z��e�]+���MZ�����?RhU��g�W�c0a�X��%�h?���]�ħ"J�ݟG�z�0�%�t�N�3s v'JE$�k��f�$�l��$F��>g�X
�p9&��!F܃T��3��V�����g C��k�[��0$���kM  ���gSO�G7r��p%�Lg�0��:���a��mN���i��&H
վ�XR�;BV�BV4<��|ی%5�4�7�,EϬ]>�� F'W'�l��'M^�z�S�i�7�玫e#��IeGnA��y��%-T��n6��緋�76Ie���
Δ�\vTo!$t��"/L�m+Y̍r�1�kQ�C4n9�L���U(4Hf~A�9{w%���]��������(�)��)4l����H_����!�e��O6�l����:)z���b�E'*��s�]M��L��e8w��/|B� ��f������|&�x0��,<*��s%�]�~R�e��8������'��P������fQL9��7R��@�4Mޑ�Pt/��\��Ā;� �#���ab�����&[J&��r�a  �<�G�v �?S ��{b 4�fU�?�VW�8��H��u�I� �S�!��k��r	6�\#�l��<�'�k��TLchO܊Joc�f���Br���UO��K��^�ܐ1ľ�h���m̮-I�:i�T��+E�ծr�0�0C��e��M-��a���x��ka�v� ��o3#��|�<�Q)���������H�Zͮo��6� �N�ܽ�X��Rf���KS+��Д=��9=A�&��C���DSU鶄�Ȑ���(�q���o׍Pd��S"h[q�;g�H������E��+�Bc�1�3SX ՠ�����-�<��c]?w���m홰v,X�&��A ����9���8V�mW""yclP�s�!3ݺM��R��<�M�Țʩ6l~c����jb.�����Rw~uLؚ�2K9��$Ze �,:dZ�+Ԫˣ4I����kr$�߮���x�5lJ�7�UU&T�,7��̇��m���?{�ٹG>98����)kf��5Gu��a2i_Ma s��I��و�*��Ӥ���{9�
l�fhz��^��!s�N�o ��&��m4����
�������2j#\��a���9���г3�H.L�t�(�㷋�"b;�KD�c��(:ʣƈ�$�K��m  ��4��(�В������:�LMXD◨=G�P3W�'e��=�MN@�'Gf��Ԝt��YJ��}�F�ȅKs��������pp���q��#~��<"M�b����Y2���p�P�r��h����Lk���+h�VQ��>L��ݦ�}�R���"*  �~Ȣ_+T\U���7殺*��dLP���@9
��[]*��}z�`GWɞ�W���)������U��%����F��S�ٯ�j�r�*o3�6c���#�d*�g�eF0�Xۼ���Ǐ�	�줎M����G�ퟸ �w�fM����X�&N�W�������l��0f�����4��Wb���/@+ۮ���p��,廼��������i�ٌ�� ���X[�Q�Z�
{�QA�i$�{�mϬ�#���^}M6L�H�o�N\�qrc7�<�؀���2Y�\ �3�����Y,�N��S%e�L�ó��$���b�{�])�{q檱��� ���"eP�1m��ȵ�Lt�q^����?�����<��C:.����ܣɴ�2�����=,��?D�����5�dnm�������#3�ϻ��,���؛�f��[o�`&�+�Z�[bƢ����F�ķ��H�
,���0q�B��{���
�C�D�6#�Eo@iv���2��)J��GЄ7�V]iS�C�� ga�"�g��
r;�D`- 8*ǻ��1�Tɉ��2���]w�l9���C��SM'��D*v��JL�d�PǳG��PE[�Kɂ֪w�!sR�us��kI1��~H��ڋJI�jw#���u��K�yT8�����Z��m���(Wמ�U�����+�B�Ƀh6�&��p�$�H��hU:�Ϋ��JT�Qr�t 8���R���	��y��D�˫_��~�^v�l�s�8��`��|��t�Z�N�����EL�A�O�[
�lrCJg�ϖGz��3�fέP�$n�7�_���Uî���C��i!cp��;F����_C��S�8�J�#�X�mۓ*i���1#��h�4z�H��n��>�<Y��IT�2\�ï�'��Y�t]����_�ޖ'�n�yA���y��{D�LY�!M#�aG��K=kHq��h��v}��#�=�Z�@뎄�$
!�f|���~(�1ɠ~��	%�!X���q��Nq"���?���Ik$�d��t�r;���>ͼ�ɋ����:����x�%w9ͦ�`����w����ɣ�ǡ�D�<�nzo��~����j ��o�J��d�G�i崇�á�sH�3-V�9W���8�����o��T��ıo�Ẍm����Hr/V,yɦUjR�����a2��t��2'$`�c��f���m@5xs1yI��Wj�v=�a�ڍA�Q���o��3LHV��������3��w#��vT(�>�Y)�`4�ǥ�F���Э������z��zy�'(-u�}%SV�Qd���217�k�8L��Y�����*�85��gm2�X�ڇ�>o6���*}XG��-��ۀ2���w��G�P�m%w5ҽ���9�՗�s�pom	�ơ4���w����.7UO �f������I�1O!J/���Db4y�|���ajq��	�����՛�l�������ؠ	�b�_�[tT �
����Kb�~�Bg�O�%)�1�)>�]8r{\���[Qx��̌�X(�I�owhP���0P�n�����yF�0D�d%��wҲ'��H/��n�|�"��y����.�P@�uZʴC��m�H���XMG���u�󰧓V�2��p�)�Y��Z@�"���u����]��N����1vv���׹NЀ����	����q:��t�֏PȨC7E%�nj�T�v2�܃�+��ݔѹ^U�2.�H�Z�e4�!^�q_�]��٤2�Q�\��#"dø:���{���?;T�j��R�t���a�i�������r�xe<|�S���ph��/.��N��,Rٙ�����qL��8��b��v�;i�����p����&�2:P�h�d���̿�g5^_@��b,kC5%aD[x�:��/}�G�����T=
R"wSK�F5��Et���q��'��*؂!�O3Yd�����<��V�>�eRktT,v����Es_S���S!�OQp�G�^�z	�d��)��p~���՜;����o�8z�@0i�b�*���:�X����}`g��u��m��
�
�9�Z�6v���>	��`)#�`�5��۷�g��[�)&,�򚜣Kz����Nt����]�׎�m��(ƀ����H�_���%M-�v�?eO��.A$�e)o����R���.��/�Kc�FH��+���U�IQ>�~�R�� 3�bd��ٕ�)'J��e��ǳy-�|\GQ`���F���q��I���P�n�O�,�!zM)+8�4Ҏ�H. ��}�n��-Z�ۙ� �8�W%�]�+#�@��8�w3�[8�y�b�f���%�=l��2�>�=MG�r�l�m��`	>�|Ʊ~-�Q�05|ŉ���|!=�1�։��ZcƮ�Zl(r���)p���M���*����ل8IC�n�έp|��^�)$�DC��FHf�oqk�D��D0�V<��qCO���Y���k�w?���2mہ���ӵm�o,��3�Pڔ L��iS��'��ށ+�X~��k�Vr�Z����<��?A��_L�t�?�/|0+{!_��]�e_��"���'�Oғ���x�M��,���QSa�V8pj�,��J���|1��L��	c��y� o5�K�Y���ή��v7u���`M+���7��lL����%*� �Jp��[+%��j?Ü�t3�>О�i+�GvG.z�kmD�@}@�+��G���I���f����1�����w�(��y�*C�g����2�s�`��\x�1%�Oǅ�������XZ��5&P.�d�A�Km���)��i.� ��r���Î{��TP�'����}=&�Z<|��|rH>Q��4���K�V�Š!(I`��"�P6)��?�E�b]����?K��cX���
b�W��BH�~���y�5ڏI^6U�ir~��.i0r^���� ����-��}�,&�`���z�i�"E` ����k��������6��ɼ�F�i7��"澒^�fFX�ڀN�f��E�����=����"8;i:JsP�A�T}Wߌ�&����i>>�sƫ*�5-Z����9�O�;�Q�����[�C53T��vo:��ZC�?a�`OM�N�is&��Vz��ݝ���avd����?��#�E���B�zJ@ L���>�H�v���[�<c	yO��yu�}�j����6�YQ���њ]D��C��<'�敿0�F�aD�F췄	���H���SblьU$�aUV�&��0������ba�%Z6S?\�!9i�J(���݅�fȜ{q��eC6�e'�~�S��x+��3(�`�s���ă����IT�:�SWH�=a�����JM�)�sY�����+�JB~K�������(�rS������¨�z�'-���d�&m���;���8yLQV:�����kz&��9x(�ls�9�P/�W!x2a���f|�>��3��j_��������9�P&V��滧�E�.[��/�r�hƶL��T�K��D�y����3r�1��#<}��-���Bb����r�1f~��'���\XH���Y�b����W���ZD�'��mG��p�����d�D�GͤG-Б��泘[�h[9�e�g����J���7M������R`:t���@/��+�N�3Q�������XM�x��`䝬��I@��z V������F7�Y�S.ig�IZ+��/o詋#en� G���4�5�o�`��܌Q!� @F�Kj�ƫ��������?��|KV��2P��ȱ������ %	1�e,k)nz���$c1 �㺵/ɯ��p�u�s��Bjϲ1��;�HZ����V+Q���Y�����Қ6Z������wq���p?)�9+(�9��86�M^���;�w8�t钁Pzv�����@ʆ��`q�6PV�#C���$͍�J\�Np�*��(Z�a����fi������7L5V]5q{\�aߑ��ش��*�4�j<`ht�����1q)ݒ��B���YM�g;gAmG�I�Q�xь�[����hz_�2{�\���RTX:)��]�6"�Ε^y�҃�7	B��J}�M9ڨ/�7�-��'�[z��m�=�^Z������V�nF������O��ug�F��31y�\��D���la3���nY/[���$~L�\0�G�p��n���kFY��� ���1d	�o�������8%�2�H�oG�<}��#��c��1�����n:*�b�� :ٙ�*��j��*���*36ٟ�0��pu/�/^�S�3��C:,��ږ[)Ӭ+x���5>�(�)���`��JX�X��~T�r�Ox�����2k���}K>s}�{8�.��QE�gQ{,�]M�..��ak���VB��T-~ �jf�)#�bJ����c�@�kA%.�O`Z�n�XՆ�>��㐥7{��?/��i�EFNŢ��غ���4ŝ2q3�j�*߿Z?��	��"�A�_���?̏ $�O<N3��ޒ�s�
@К#�p[vi61ihٙ���RՈu|�\A�5��\��$�K�(��e���~�K6&�p�F����?a�F�B�O.��N�5���A��ކޤ�A�J�Ut�-E��{0�c+��M�K�GQ��u���O��ե���ʄi�d�I	��2Y�]]��N�!�$~����V� n�Pd�<��{��4`@~s�<Tl�U�d��I;ϵ�X�j$3.Xͮ�`�f�����n#ݐ�o�W�|`��&��4�-���/�y�fCmB���iν�7�ђL��@���&�F���h�'b�� ����~�;i��6uI���goH�����s����N���1<a9�����{BLOۼ#P��h���!>��N��ر��U)���}��\�ǯS̸ �B�A\ѿ��ѝ�W݁C���4��w[��Gs��N�9��.���	\�N�Ў�0i�����b�*wƢ��µ߇�z�FJ�v>�St��,[��a��w<���n�b��Hӝ�ų����$�}0'ju�Ή��}� �6�f��w�;��lVS��p�*��s�dG��f�?�Ix/a��*�~��%|e�X,Q��{�f�B���8笠_�ֿ�@t��-�ؔ�i�C,��.��[�����h��C��^n6�-'�
'���K�l�i�41R�HV��إ+G.�f����Ռd1I_�Ԫ�n�2ֲ�9��L`T��}��eR��+iL�`Z��	"�c��m2����jWM�ҷH�y���� B���������������>�D��|)�ٳa��P3�f�<������|nN1�� J�6�L�,�_!��XI�Jp�i��s:�b{Ģx%8�N�a��z �s�r��6���h�Cb�ՊGg��y��Aq~W�{B�Z�ⷜ���b�L��8^���a�1r$��q�c�MW�M֓Bn�Q_+ɖ�s��]l ]L��?7G>rs�(���T�E-��b��޸�d�a�A�[�p����u�|�AW�*��o�ͯ˳3"�-�L����)�"BK�&+V�E�U`��V�dQ��>g��JԵ8%>M�]ڥʞ�l�"�ż[r��]��F��O�6ns�LQp�T2��o�|�Paԇy`m�-��b���l�O ��,�Q�:����n`�ᦣ8�����0��i.�ݍ�����]%��D����oʖek�+ [�(Ow�G.�j����P�p�/�ckj��V�n}����y2��[L�Svj�i�Xв=�oin}�W����)c$�S�n� E��"P7���N"/p������1�O�|y��z笄�6��B��*íX�:����R�����F�#T�lʾ�V����ݫ�T�{�>���(8M-%4`���}+��6X<�A���>k�@�JN�����>&1!qT�V��R�t؝�`�Y��>�U|5�uAV��Q�\x�Rh��v)�H��ә����x6^(��9�G�&֘� Ү:���N.��.��&/��* ����J-U�� `g�qo�oO�\���ZCFm��vT���Vg@�h[�6�D&���]㒙�C=���������K߃j%��6�+���A�ܤb��}���T���7ce	_��E��2�<+�9���OŌqP��X?���%l���N�Һ|^Pb�<�2ku��gR�+�f8�|+�/�|��5;7!CÜ�Qhy,Ccg'�|�0�v�b/�R؄͗w��Fo��՜�:^Mi�E.���p��������b�*ke#���oiJ���)�}��)�ab�~0�t'���[N3W{�=:��ў��������y�G��V{�l��_��Ȥ�.�(^j���<]�xV2
�u�J�蒍�%Ƨ�aLk�ؚD���/uU�z���q��N��WP��/��'#���G���f� 69kl�<�Ta?>	j�{U/уm����'�>�Z�E��ܷq�6�:��h�Md�q"	�c`S�	=$��z��u9�`�o��w!����\�r^���<j�q�9w��R�ǖR��G= �Z���;Չ��w��}��Kx�Nta����MT{����n)I^ʑ�Yy�#V����D�d��J;w��z�b��Y�����cI@�ß���ː��3�-oZ�:X:�(���y)�qJ�6�a��s�^����8�zM:;���F���\��;6M4��^���1��X,��j�W��A�E=u̴9#L��s�;�<F����ud'ǔ;١�9 cN�DY?��h��#�;�+K�F7|h8F��Y�J��!G��]�߫8vn���(\7���� �������:C��|���v��#i	�F�~�㴛�&ഏ��ߊJ�/-Ђ�b�Lt��)[I뙩�x�2�֦Z�f+�_�-r����b�|�`5��ù:�m�(�fvJ>rW3�sW��m�`L|f9���65�L	A-A@LIM5��7�k�}�[)�~���n:���ǚf��A��w@�T��䟢	Cև=cҠ3Yɇ�!�0�%'q��\��Qo���e�c?��mTGꏾ��8�.����6�(y���x�ǥ�GȽQ���A��k"7z44�b{��X������SKqz{�zG�E�qUmN���˱;ƐS�a���C�#�:��à�E���6}�������^��g�^�_!KКŘ���GX*�cN0M�˫zcX����OU�ޡ���1=�\�'w��|��O �����y�Y~��ɣG�WS6��#�RP�Ar����A�;
�)W��N�M��#mM$�������3A�M��bO��$=�y�	���L����9�څ�S��A@/^�T��[@C[�1�5@l�#0�W�����ò;Xv����7�{�J>b��*E��T�L�-��m�8�񨥸��@�51�Tq}o؃)����`<y�P,e�8��8֓ Gc���[�nLu��?���G����ݫy$�˲�D���LJ]V$�J��jھ��i=^��7<�M6q���� 3&@̶
����p����@��.y�JU�,YdT����������=�d����G�^���'��:��`+V��iy����m��"���B���^�_(}&�#�9���|�'�Bn�_!yu󗭝�F0u.A6�*}N����茋 ������;hfEt:+h`㊡P*��U]J��������_��a�M�w�c+Y-�x(�\_^�e�R88uѻ���Nt�/�5�(̈Ӹ�Ũ��@w��ހ�#���T|�P����u��o^��?��i�Ƙ���r����ˢ%/�0��Q@��E��z�[��M�H��}J+n���ٖu���
��^֭,����͕Y�(c�z#���1�����䃆�r����N�6#d�[�_X��O�5���͞z�>�ϣ�N"�/ D��8�*��
b	�����y5֍��*r:��#�L�f��htkU�l��z����ǋP�\�������=�}iG��C�U���u}#��9��o��Q:��3�1��5>W��=�E�|	:�
�.�[�.��C*K�6a'f�l�m���.a&q0ar��,��h?��氿����ts���������?v��g���;�(�խ|������L��1�.�����.��[����Bҫ)2]'Z��Y�����X�KXkd�����Fn� �ơ%�J�i�؀���O�m�����s����V��˖�U0n�=~{�I,����yBS��daA�pF������Tv�"?)R�q�l�}�2n0�n�tz�+���/� ^C�t\��@[��ȩ��Q��
>f"�F�g౿k��r��!���+o�Db����9S:�`n���85c$l�"�-Xl�h�˄s�%�%P�
�aL p�6	PJ����,z�W�߃c��Ym�c�p�&
��7b�{w_�ۈ��&1~M��[

>4v:�H�6N�w. �vk���ӫ����@7���!}�8(��R����'x(��ԄY�K	)@c�/ƹ���mZϐ�4�h���<��z�X{����� Y��"r:���r�^IPjC�D���萵��Hw#� �lԿ���X.�v��P}�P���BY��D��N�� UM���1�e�H�]ʝ�ZԎl��"㿶?���_����2����#
��f�O���2�����b��,�n�s*
F'A�SK�sy����EWN,
E�Yt�&�܏������Bw�7����Ӭw�
q} ��ೆ��m������(w9��V�K*9s���vp� ̌(�g�6��;���ԐS�,�{�l04��Q\��x�#c��v\��s�ʝq",^�ĭ:;L���]�7i�O��D�LT�O�m����Ȣk47�����/�9gf��]��<�P�^9�<%�r�+`����N�����	͋����b��ڏ���"C��$ؔp�����F_t�e+�Q�ݚ�|�ϧ>o����C�x}�	/����Ln;�%�@uWp̕�5-�`��������H..w�j$����]�*�x�����ө�����z�]sE�Oư���1tܬ���m'O�����F�{C�uGwZ+��j$)����JB9�$=�%L+����t�,�HʈY>�qe��I���5�܃��*u���T�$kЎw���/�����\tvC�k>CH�"���i�QC����z�ìvn�è����T|�;w�+��jǤ�z����E���uh�b����?K���eI�G�/����%`��e�_/#^�Q�����E�1���l�?R�����O7������-��S�y���(PA�/p�I��*��O��VB�<(h�7�YJ��d��+���_B��P����B��TcC5�{�z��#��9���Y�2��at�i>�����UB}Y��b�#e>�rI�/lX�BD)'4ز�6��԰�~���<���J��˝��t
XW��^`���V�*��Ǻ��K�m>.�?��l�j��!�x9۝��:��`��Q`����y�a�[Ű��~���`Q~T�H'/���\Z���Zf��sXb�
��irܶg�p
����*��ut��p��'=a?k�]A�����A�*u���Q-��hn:�&� @6�İ�W��߄ԄZ�^�		Ǻ�A��?n���A�jUzo�Y<$��N���懞�5����.�B����&�%�箢��M�*�5��׺�pUl{�����ohaGPx��	3g�Rڮ����]�B ��I�BJ���ڧ���k���5����x]	�E-�>�� _M�۟P{[���:�\�Z��U��G?�C���o:��U5V'�����E�V��g1������m��I.^�������4�4�<x0}��3 ��
���үc_*{���r��DWKYD���SOX�SŪ��"
��w�D���)Mi�[���3F3�gE���/G�NM����8nZAn��R�s�C�"I�0u&�aA)tX�р��!��R-HVT����L�'�,��c�S~�ᆰA�9��3�%�0bs����a���҉�\LҴ���Jn��+5oS���ݚ�AB�����F�J�D�;�?�d&-�o3�ʵ�j�R/���{�a$t�������6r�v0��X��)a���x;|�!�:iq@�%��1�o��;
K������W�xE�r+6uI{��ih�z^��^"O0"#�.Sn k�2.|pҲ�S}5�Q�?�/����&~?x���.3���,c0vN�-4|�O΍�;9�_��� �BQ��R��qQ�Rn:���k_Xa�&�2 L����đ5<�417��u9:��I�Q�����{fH��x,-�A��I��/�į���>�V�ɈQ�n
6P��`�b�.v�Kϊ�ި�b�+�
�W|�0YQ���\���)��;��fz��*)��G��eUC�����Ii�V�'U僷��x�Sn2[��]>=�����D/؛��TD	��IE{��7�t�u���o;տv�ZWT�T �27��wH`�EW�ؑ%'5�BKޜ=�"W�(O�@|u�����),���}~kf@>	ZMq�!���J���I����N��
��'I���&^��	W�e]�|g:��.����p��<�������`\#���{yЛ�c�4�G_a�LQ��>��&q��;}`7"���.$)_�ؓ��,���t�����G�M����9�2�V�+���c֮�%���'[���� �g��w�VT��j��d���{l�u�5r5�pd*Z�Fn[����'/z��S��er	��$���A�X��ā�\�ɮ5��/N���ApT�%@����:N�(�����d��>}[�����	t�5�B:�)�2���:��S�ͻ;�2d��11��1����lW�Vo��ap��ݷV �g�E�b��$�� 6��'Ǽ7����+á-'(�?!?4UJ1�K�d?�Rs��GU>@��y�|OE�{�-�.kJq�MI@�(��@e�]6�X��g|�F���-����֮�Jp�)W^I�5F>w}�F�;�L�Y�Q)�u�c&^0�FQ ��(��8<���"�Z3%-���97�����SM�Sա���vN�^*�9�=���np����?U����wj�رvҢYY�ހV�wշ�}�u��!���"��U��i�)�
a-y��7su$�,C�����K���ԼxԹ��WK��3וeya�����?T��z��g�^~���n=}/��r������R�Q�D��-We��[C&�N��.2?׭�c�e��~��wլ~
-�	�d��װ6��8�����,S-nM��6�K���.�s�����;I�.��5�'L��G�|�,I,�wh�[����=�m>i��$��?��5��㷩yZ����$7���]�ѓF�<R<@��1��!�����zc���%�v���F�k����N�R�y���{H�־�y����nѳӇ��8��W��ƫTcb�CncB"1���2Su=����>E<�Q+��(���������^�C��O#� ^w�i���g�Of�l ݄��6�9 �����=w��~#�MAE�b�@�^j_�QD����>���'PO�P�넬�
,Q����Gv��L�(��$������wݛOO�K;&|��S���]�t�.nL�Â���V��?��`�JO7��	,l_�3mE���_5�\&g�\�[��.
��ü���g;���$'�?�=:�j]�F�o��AG�0����z^}mE��D����Ő��7�Ưvw��|���N�̧τ/c<V�YX�����K��������2�7�?�ES"P21�<����]��s8���I�*ғ�;V�1���x>w�:2R�k-�vNt���WVO�h0DXE�_��Hс�����l�{�ir��ns��鬔G7�0��8ly��4�"n�%��E�����b��)w"y���݌�J4|�֟���Z1���;z|�5]necT�@�t�g��	�=e�Ȭ�6�+�|+S���x5�������M��ց���� �L&%�Eڼ���OWbC�5d��J �d�3����y�ǧ�ܩ��]��7JUyj�{�LRc�rGr���'9���6�:R�U��V�뢦9]R�?CeQ�n�T��J�t��
�\ŗ839�ܧhnbI�x~[� ������5���rq��u��s�H;
���ڲEKC�J��:D=V�!L�j2mY��jB�'����0�G�?j�b��^��D���5Z�����,0�;�m��_�6��~��A6נ�G�*S���8ڈQ>uG�ڡ6$��/>�Te��{���l�_��\ɡs�WJ�aǧ���@�.�c/�?�4�� ���s�ǻ��O��uy���ɑevNM�pb�	'>�'+P�
9�_�聊l-{Z-���]��/9���ef;�7|���������3$)����C�l]I��O���m�j��H����.��:���
ћ���S�$���h�
�)ZhdV����x��4ғ.�vw���C~�2P<$zʲ0r��[&�+�^jV#�^��k�$�1��Ӏ�¬|��ԙ%������-&#Q�;����,+i.��x�-����D�_Ւ��cQt
O�/���� ��,T�~5~C:��z�8���3%�5$k��h��Y�����#hֱ����Mp���q#5����k-D���D]B�ؓ��qL�P.Y<- XI������$�;��2�U�`>γ�·�A�&I>p\�?�V���d�} �G.����L'�E��ITD��sN4'W��>�uyM����kcvo�`	�#�^L��g��SW��ȡQ�v�Dd�	�<gm�P�=Gp2	(������Ҵ�М�r���xl
9��h1�
�B��1-�e�����|��縸���}&�T�?i�RD9h�,#��h�rq����K+	ף�F/J1G��ݷ0�w�,�>��J�Y����0�F6l�M|=yUg���^ �C����'�Y�}�0@��CD�w-)o䐨F;d���|�
E)@6��N!��N��Iq5pԗ��~{��^�
Q;`CYzz(_�Oў�����mÆ���.d�u ׾RG��@���E�����r��Q�q��a�?�p+��t��(<O.��N@t�4�0\$�M|F���������ϳ��'��0��P�L~1ey�ƂUl��6�MPs�l�m�>Z;}Q�OHx�hvx�)������7
����0�Fֿ9#z�yH��}�*�6�(A���#G���,�xk���x�N����'o� 0��G O�J�X�S1�tB�u��R;bT 3��b}R+�gW���t� �'̈́յ�7�!� `#��p|��_�r'l�5)�"ַhO؅�s?rP�`睏�W����4�m�iw4��^g..�4f��f�*h�ye]��^^1���OjR�/���=�ҭV�of�	L�0fO~�l�L�kg�x$`��x%85*�Ұ��/���JU���P����%��a��Y�f_���p�8��	��c��U1W�<V�y>aEk�ɸ��Z�����gK}��a�$�\D�]�$�Y��jb(]ښ��9�Z= �U.T�^���פo��� �uPq��oE���|��-	=H*��,p�G6�'�b0��Q�?b�V�骲�����Q'��j��c�qű�܈�ri�!3����)Ï��,視��}�g������������c�ŋW����A��������F��cR�h�q�ד�(Qɘ~YGs�b��<��1�{(RKb�<����4��l���*�G�
�]	�Y�F	���L4E����l�� ��6�G�8O"aX����}Ƽ�h"{��:�5_��c,�9S���z�dҤ]ҙ� �\�j	2\'^�!u+�������8��V�2��q��d�3NHsr ZZ�E��*�e��y`#���]�<NH*�������P>CK�'M���N�S�D��|�>��lT����H�.�F3+�4���R��NX*	ۉ����8�Ng�A�?�#��C8h'�.!����s�=�!	��y��e��G�V`���y�md9�Q�SZ%l4D�%�3�?��<�2��˞<7FKר}��v�,��=<'n�0��-4��ܫF���5bXr�r�QD���=����`$�����\+��$�����������g��>1�i���a=��v��Rؓ#�`-� >)~ޥr�{T�%!�Y�����n�#�d␏��+��#3��m�Ȃ��}�^�*ݼ���A�=�1h�A"/��k�����Ds��O޶�p�~ gk�stae|���Fn�tl�АV�>�?����9��#��Ǣ6y�D��^�:��P��M��b�k~��v�8���Z'�_W �L��1�~��`?�΢��?5����~�x�F��|L���ᙵn�G�n�[.�Ki-��*��5�){���G!杏��B�7FA�$"�SEA�S��g��w��N�-Ը'yn�~��5��ۏ_Ћ�K5p���j�&�__��C��*��\"ئ���dI���Hc�k���Ж |S$2d��%f�����s@6m���=|]a4ڰ���?�권 ������Y�G݆��,~?��ӆ����� �6��m�S�Ծj��}D������eD��\�C�/�VA���Uˠ�)f�'<l����Z������sH��<f��.v:dp�χ��.<$��i�<����l]Z�X"}W�����o��xi&�2U�"3�6@a�6h)a� 9'>U�:���H�KF�� U�ɮ�����G�w{?u�=�=�5g��O�9*��q�} _�{H���f�I\�w�&��֨`�ZAe�����r��^�u`j�W�G{� ����8�-�jt�0�)�p.���#�Hך�4Gp�w_�hX��q�I�ݠb��;�ɚ��A]	�\�L��)ɨ�!�l�D_,#���vK*^7�JG��ھ�c���=����[lIP1�?�\TƢ($;��̞s�J#�����`>x_�<_��Ĉ>~ p���G<���@��V�;�,���O�GdU}|!)����a��R�2�b����H�1)B�q�m�����v�nj�88:x0�ݵ�7�Dci�ld��!�	l����{w���5b�)���r�)�܆�����6�uW��UyAl��l<��M;˲-�<�z���|��Y]F�DZ[YS��96�G�����t�_:�O�����Rr:�HK9b\�v-���J~������B���~P�C�,T$"���9��@8��-z�E�bj��ߒ��ͫ���,�ӈ�O{~͝/F���d�:xw��˂�%oH��3 t69��� -�LsJ9}-y���SA2���5+�~RT(����U��j�zM]�C�&��&<��R'��b(�Z�����?��!�E~HK���M���7gan�m�a���{	%S	���K����/}6[Lv�s��Z��H�0��D�`oP�����֢��^~���&6���� 5�W�L�N��]�������558�����Sz:>��(nXԁF�k���~�KZY@�O[��C��Sc,a:]�ݤ+�]�M����='�p�W�5�H�{�&}US��) r4v����.�`��U���K0=� ��&Zi�9�I��@�@�,��:�����B�k�=
�i�U���<�P*��[@Q����p4U�-�Ț/�iUy��܅8LN���n���
�3U����vv�^���b�aO��-xv���g
[��K~�b��=U%-�#>��}1�r ���]~���hQ 8hQ��{'Jhi���IoZjgɱx�2���gE�j�˗�ż�'����aN�'N�n	�*uiSA�\k�y��`a'%T���q��M�'���81��i�5}����t���w�8b��XFw�6)t;��81V�'7w���f��ˮw��X
�N�~�Q訵��F|#�V�)�L���2��0��Xަi$��I>X�����Ւ`N��'A���ALV��������}O&�)�����Q�z�X�%<�l�h����M0�.i��lM#�j��G����Z�N�0f�RO{�;�w��Y�3|�yY�L��X׶���ĘpIX�-����6��ʤ�y�4��xv�IH`:2w5n&��qyT��n���q�����w�'{&M���r�l	�+����d�x��h���fd}0�K��vY1L�Գ��xu4�T���g��%b��/���3�[�	�$��y����wF�~��;!�ɖ�}�$��H�
��hʱ�U�=��)8A}�{	�C��F��]�N���&T�_��t�����&��L�ֿ����V�Y	Q�Q�+�J��gj�Z�?	є���5Gw�Q���/X�AM���ϫߢ)E���o����\����0ɈL!�KK7�5��{*�Gk���A��.�lFm?
��
[7"-�!���ȣ�-�o����U��(`�����.�'������.z��6�5;F�̣�T�y:��A�����=��zJ<����������@z�E~�`$c��7���b�)�\��>Ќ�lZ&O9a+v��`��*����<�(e���r�z-Xu�j� :��b�EZ�v��&��'�0$m�@A�p��Fv�a���ԙ�Q�A컼:�Q��~:	�!�7�z;�]#3�lT\���s���+��C��b�]s%~w]�nS�o��:}/�]��B�	
V_38e��&�=^��S����#��@~R0Ґƒ�0%}� �ɺ�q{Dr�f�7��� �P���}"8�!f��8���<ٻ�����"�Ӏw�rl٬�ܓ�Eh q*'HϐMp��P{ʇ�\�L�#�#af�a �_7O?y�������~�\��g8-�Ra㲳�����g՘�bv]L�)�b�~��s���e��J_��'o.�-YLZ8�>c��0V�,cW��M�����9�4"|_��W3��Q�0�O��f���LZ�r�˟���id��cҧ����ɲ�bV���⃅����g?�T�%!�D���`�K��z���Z����W�$�����!
$k�/r-���o{�pu=x�^e5���Z�vH2���b=CL���h|U�2���,��k	*�j7^��4Y�l�����؀�3���*�F������P�A��,-��z�uQVSo���fY��U�M�Q̍��JȜZM~r����ъ�i��og��i����.^�����x��R��������6������S ���c�3�%�Q�b
oNt��-�X��;/	-/c��i��7i��Tx�4��&%󀊒ermPı'@N1VY�f����1%�;7я^�/S�g�c�v��+�!"k�������U����s��&����^yxGJM��㴐j��ү/g-E��xu|�[���m��r�9?Ôn��I�tJ'a�����ے�-�S���u/Ui�~������u����B�B$����+8���uLy���e��F9�[p�E]]��iXkVg� >�F������������;a}�7�3��0���q*^/%�����%���n��P�bt�l�w�(��T.e�XK���H��Q~�n�ÃPXY�HWԪ'��s�{����_�H-aG����t΄'Ma���#��xe�J���g�6��� \<%8q�[A3"������w����2�!>z��?+�o�rNk�����nK�9��o�څ��m�!�R'�	#�Gj4s.z�B ~�j�j�Q�<./�"��+1�7*��$?���6L��mE�QL����ѐ�6{��`��O�	�9'3 %�l���eƲ��e!×UP�	����Z�"�o�`jfnr�Q�V.�՝��֊E*�fP�����m~���l��ș�ը�L�̷D��U��7���}ER�m��W?g�J�M��BS�P!Yׅ�� g�(������/])�9{]F�w���Ϝ2,V��vn)�>l�rV�_s�\��]V��㓻vhKK<��	�eh����<�f6�yf@?&]�S�g:l��]�ҳϢ��L��-���.�v����X�a��4O�/K���1�Y��k��a;����.B}S 3��ݦ��w5��G�
������r�K9�:1pp������|�GX���U�Ӓb���j|����/�J�F逶Q�!�����J�J�SKv*�.8!"o�����O����9A��B�f��@�u5�Szֆ��A�|�ؐ��_B���	6_x
8�vU&����P����k��Y��#�
��i�\}R��q,���ע&��1b%$я?P�Q�-s,s��ne�lJ4N��ku�����M�����4�(S�?H��y�cT�jma���Z�}�U8���|�Kl;дp�}}г�lhT����U�,��8������P�ml��{f���?\c!=|A�vF&��xm����>V���o�%���.*um5K�D�z�����qE���{=�.��z�%Z!�@����_X��X�-�)�1��M�X!�+1��ί #�pQB?H�qo���s�< ���3�$M��]f�[��<��Y��]/�����Fx�xbbf��ֻ3*F��o�Ք��iY
S��	�8ֹ�A�'�6�I��-~�cb=�#�D3a��)����9�D��.��̈́i��[ϹV�����q0�p�-��4W��v" ����nXgg�,=�4�@U��I[�c�
���6Y)�:i8�¿$���]�<ܓAQ�WK�2�F٢F��T����h���E��o��ƍtav�����
/�x�Rf��x��c���5�Fl��;�g�d������n�)!�Gނ���|��MDkU�$*,�p��ًگ^ѯm�GV��u�v���}�Y�e?����s�İ����Z3� �t�W�>��P4�aq!�t��}�f�� ~��n��󽌆�@d���<r��/`���$o���XC�VZ{�r��b'�ꯅ��Cf-�Y�6 7+"򽷩a�^� �l���I�Zf����+�� �ݴ��;��p�(=�%b[.���#��Q1}qq���)��*�'N�x�b��/��5-ԝq3�%�\9K&7@ŘA�:��bb��ΐP�֓��c,��G�3h ��c*f֥�U�â�Q�ܵ��J�ϯ10���q(w�?.�	q�6�ԗXv�������x�T��\�j��BK�F��<�<W��HBl�^���<\!q� �=�ѕP�+���G����0�����\9Ѽ;C1����E�F�>��Wo����ٓ+^G�F�TaH�j܆n���0cY��mn���˙�qq}Nid{���6{c:�˳<vɷӮ#02xL���#5��@:�,m�z���>�CM�_��p��שf��H�p�T�X ���>�a���j((�pV�~ƪd_�K�LgL����.�dԺѯ~7*��CF|�㐐P�E���������ڶ�#E#� 8T�x;�oLK|Kiٜ90�^/6V��/���ڊ��A�c�Q����ZG
��r"OMR�s#3��6C�����0�+P���̘�M%�ٹ�d�HjH���([�!����vtR+���7D2@;���L�o?3pD<��C	19�S�oYv1M:F�uqS��C�M�VS%��Ӛ6�����Nb��q�͜��3�l�٤j��߲?{��7����*I�<��T�5 %,<���#���T(�M��O�i��%Ft��q�U.�KL��Rh�ٌ����Mp�iM�wd�fsID̨� �����z��c�m�:��L��SQ����o�y�KQ�|S#���u���`MT�^~q��|���H`m�Iq}�=k^�����ޜ�06�3�=�g;/)��[�n�*/yx#eQ,Ӄ�ݨx>=8Ћ<ď|��Y��i���m4�
gk�d.i���X�������9Ќ,V�+�>�8Q^FE\,�>Tg���O`�-���%���)H/���F X��DNpZ����8����l?>��'����
pS�lh���9z@��66K0�DQ�$S�=ȕOA�}g ��Q�?d-�&���O�Ka��b��N$^�a`��Ý��շ(
pP��h��>�y�;1"�8X���8բ(�f�}�b�s��%G����b�܄������F0�ar���3>�FޯQ��C��@�VØ��&Po��q���D�v�yL;�O�q^"��R{���S�!�ly �S��&�aǆ޳��q��#�l�ǟ�%P ��<�К|@���T�F6C�Q�?/;�'�;�XR�s�]hm�T�[{��I�?�R��|�9���ܟ��8�������h}����ӭ����{=o��(���m-�j���9{L^_���V��ZL�s�MPC��%ز��*�,��#��QI�x��?P��&���i�g"����O�@�?=_��iNk����jii�φ�R-'.�vOO�3�w��\Z��S��19�%��x7���
�ء�`!�J}}�A����
��u�FF1 �L'q��=�S��C�jߺ9�-�X��.S쇶;��Q����3��U�2����+B+�0J��� �@��'@����/�/c�kS`mˤ�rb�*�P9L�Ƣ���u��:�=����\��X2L �h������k���_i�J������u������^#���k�3!�j5�p��q#�1i�Ι�(�ÌT0iJ���?Y� �Z��dbv�t;�Z�ί��2*�X�'P��T�~��R�aL�9!� ԏ�:�P�)�����n9�O��*
y̘2���F��
��5�Y��R�d[fta���2�[�|�IX̲r��Ŕ����ɿ2F-��mZ��GV0�GH�X�m�+�,'�h'!v�&$J���U�J�d��2��5��Z�(!�j����)wlщB�q;I�=�#����*������n�sW�����K�V9]p$��?�;\Nۋ��9�x�T']�ʮS��B�{�ث_�5�ݫB����G(��w'��Ѹ��I�0�Q��^���rD	HZ����C�y��>�r�g���VW�(�+�_I ~�����7�n�e�������,���"�$e�?���̤�n�h"��/���6|3u��[�%ʡqb?��-���/)�W�q�q]'��Y��̲D+�g���F����r�i`.�#<�8xW�v�e���3�ďbW��.�֫}�l�@D�1�^�'��a�B�o���s��d,*+>�˙Ɍ�g����+�˒���7	@��8�\�<�".hH��b�Y�:+�J�z<i��Y��Y�)�V��c��v>�]��D1���¥����(�`E���=��̕ )}�1C���}a��ͦHBǘb��9f=cl�J������^h���QG��m�V��E��CjB����!�Ro3�3�P$󜥇����j_�����a�ǰ�#ka⏹D��6��I�p�cQ��|�U/a(l��:�\�䮆���㲐�[�?gBS;�[Z�	���7 �lQ���@Ξ���>t����#+��4#5+y����cG�)�V����Tm��^1�����<�Z���R�M�'
��1��G��ۚ	}����*J��Mh1qqs��l��i�����Oܕ�*N^a���
W������$������������.���s�ǗҾ4���z��גq�gR�';-]� %�Z���|}��nP�5���m��W��	���m����%2�!3�-Z- �ى�G��G�|9ǐ�#��\y��_-��E!��5m#�n���'���� �RB�]5�;�&;���6#2Т���ؐs'L��d�q�����x8'�]n�S7�</73�2w��yeE#�}�JM>����|�{;���k��ά����^�=��O���Nߐ�b<#���t���>t)��Mr��,o���YЧ5�L[eI�Z�8���^۫wC�I$�H��#���2w"��JQP�|�&�)���G)4�1+r�'����ב7 ǈ�`�����u�3��n�]}�>��-�*�x���v?,��-_�^�T�E�U�c���A5�o�`���;�N?�#g��=,�j�����Z��M&�"&�$�^�JaqPGa����KӪ_�G����I�46
c�� �P�=��Xf��}�l�J����Ϙ߯�����N<��sBd�T @���:b:��Y�F�`պF�x�t7������2������3�g�����̨?3���-^���P���9*Yb�l�z\R��,z�m@Zu�,����D����ݧ����j���s/���B�o�T�J{���١HP�TxC��"措�q�ÂԊ�h���U�
����]���Њ���
���BoIS<=YM��s�4N�� IT6-�`Q�f��{/�LRnz����'mR�����c�(Ѭ��	���g+�lJK�i��0V��a�% /��܀��v�D��y3$嗚�JMF�@�8���^�q��o���;^��F�x����B�X�h'�*XB��㫐����5J���I�
E�N�l����0���m�?W��F�D�F�yR�=}#�XJD�5�F��a�U�\��덲�?���M��ܳ�ٽ�ډX�+"~x��t!�����L�v�{<� �i�9A4���[`��L�V�	}�)54t��������egJ �x��k��X�ijO ��E�3Jb=$��a���;�e�o!�D+Fx�&���^���G�;��D
�6{��ڹ�=����aN�_k7���!�p��޹�it����C�X��o^�n9�?��a����0o�c�$Lݖ��65+%eoQ߈����A�Df���5�mJx����װ��CU{ �����hn�0�(�I�
�b�(�	�$��ފ&���������A��pC�Z2�t+E�x��1�� �h�չ�w�����H^�G���ĪUWg-���4�-�����|7��x計Rg�OM��6��P�K�w�u�겣����{ש�K�@���^�+a�V(���*z����4r���́�`:�_��)`X����R���˝��%tPA>8��Oh�˓�w��HC�isu���&w\���[��̧�9�hE�dϐW��g!�V�EK�u qN�D�<�i�ζ������EUM����=\舉*�N��Dq��Ьr9�2�z3�;Χ?�:r�^b�����c�:��+P	'
�[�:�e�������&EJ�FN�����
��!�
��].{N�6�	aL�\�G1�
d�;����x�x��d)����N\��u�H�T�yO3�˝D_F����Un҄��N�(Z��]ƪ��uv�A�DZp�ir1y��+I;qM�ܓ���m��߽�t[a>Ʌp�'ё��}s��4/lW��Q��/�{9g��)2�'E������ɒ��LA��DxI1+�����A�	��	ުq7�G���f�`ۊ�-'9Ma�S� �-��P%����T����$�Gf��X���[�ڭb� �51�:>륿�f* ���S�Ry�,n:z��\JV��:�F�a��	p��q=	�D��H�B����y㫽�����ջR ߄�Ȋ�̦�,$L��:*�i㖈\gh�5N�ᕃH"��k��
0@)��wd��{���=��N]���<m��93���7H?������S�%6"�	pa	̳���F�ȘI�+��7c�?��^U�����.�����פo�Z���`�q�DA�#�d�-����3���t���&$N�����5q���br�`�O�K4.\��3]�S��0�F4ֳ��%iN3�Z�=�_-�f�l��d�/�m/Z8�"lv����Y"#�ȶN���Z��n1mlȀ+��D��Dk�C:�!�msͲ�z9�sie"F	�$��3a���]�o"a�O�-)�/,s-�P�!�o�o��瓘v11l�L��͡�@��u�)o�٩c	�;��,/?���۸�Z���֝����#>��W��I)�Z��|s��/�G��NX��^"�5�Q���>�핟����YguB���ؐ�g��9����������,*-9�s>�ӓKDwP�:��tX_쳥����jR�%��mΊa�V��]�,AR�l�3*=���ʭ|"FyĈ���=q_ \�<��t��W���v�Ȍ�6�f21kt�+4��6V{3ϣxo�̔Gf��1���<R�c�wN���ǔ<���*��1o�=���d!;�k��6�D[)�L~�<��B�[��}���A�$}��'�c��4��_�Iz ����>�>WN�;t�0ho=ھ��x����G��@x?�B�~S_OW�2�I2�����ۅ-�"�*������k��?)�q�q;+�h��O���nP��H[��k�u
Bw[��X���w����\��[ �(�^��C�>���ΐ��f�C�\F0)g��̩YeeО��ĳ���'��QR
`����"�,�tjJe�uv�c��b��&`�?�S�T]�9��#Ձ�Ú�/J�%u|��N*�r�ωgG Č��ғ����3z���	:쾆°��j@�*���]X��D� Ŷ?�ڶ�y�"�p�����S4 [[�no;T�l'`����P�Hn�;8 ?�̏S=@��Ԫ{�}��͹�e��n�SR���e����\�ш�� ��JZˍr������-O�\l@���G?�#���K��"�\o�j��c�:G�./�}��"
�`f��mk$�P3 d�&H�s.�~�`U�?�ZG��3п�!�7���@�&���]����5����[�uWG�,�S�Q�,��Y�!]-{���e>|k_�k���*��ڜ۸
��7Ea����ZeX�$��wi�l
�c-j�T��Q�VB�,��=?}���Ɲ²�D�py��V�����/���)���m8s9^�2�h��t<zd�IїI+!��􁗏��?���K��c}��n�m����U�ש�� kTЃQ�:	����|�)��(��\Ԅ]����n�7aѓ�LQ�c�*g8L����Ssi�N�W���D�ԥ�ޛ��Gر��6]��<�ٳ� �r]X�܏�b'�U�ɡe��$E�s�uI%�+7�DYF\	�[B+�Y��=��ذ/�ۃɆ��z��^'���t����~X�/2ח�hRfPX���|���6�_�m�s%�V��!&l��ZY�Z��s#��*=B�=O�2mRH�A�ȩ+W��W}.A��c�!��D��y�36a�m��\3d|*dx�!�b45� 7 ø4�aj�e ��w�;�^�Kl}�d��l@ x��d��?t��SR9]�UW���6�Ӻ�y�lU�?�e�
p�Kc�G��;{K����5�3���ih��U���(�58��̥WJ8}ʠ�![Y:[�Hy̭����(�Ŵ%��zhu�$��_�q�9!V���z�	�����sx���# �.�PE�0��2fI��p)��la�vD{Kf���<��HjFh��]���>K���ۣ:!����y|ɣ��9g zg����dx�V��-�8g�"o�nZ���UО�S˕��P���[�=!�3�9�(5����TE*<F�+�h���ţN!O#�Ux�@J�`q�� ��Kg%[b?�óF�&[��)M������g'��~%��Qp4����z�
��>Gt�y9�7*1]J�M{4�b�M�x-rę��y�ҁR�ɣbh��V��Z��P�?��i]X]�.��2��BM����q�L�N�a5oI!�I�*6[��T�֧Sz����M���bB ����߬!e(�2* �vT��r�Z�h�Amy��ނ0po�Q*�3�P�o�Sj�0���d� 6[K���瓫���J��H�J'K[D��V��x��f�7�!7j�@��|;���J�w"Tǝ�����F�����{��4�aP� �f
S�x��C��j���T����z9��簶
�b�b]u�3�m�?�R��O<h�� ��rNM�B�ִ��|"��!]��>2��	Fgl����#ȱy���[���tu����SY���Umyf�լ�k�L�,k�����q�o������Tib���(�R-@��]�*M���	:�����	l�ff<u"uP�5j�K\��f"�]p3,m�k�@F��h��d�'T��t���9{��e�J\׺���0Ǜ��D �9�b��A�/���v���3�ֆxQ�(R�ܭ���D�a8����M��C���ΖR�?�{���E�.���izS�|����*��$�m���?Z��HQ�]@k`�7��[��Ko�����lU�`lY�n���l���|���V� ���忇���5g��_tnX+�`��Q��fM�d)\�TL�	�N���U�ݕ6�:���	�@��4	ۮ�5�i@��H4��4��G*���8)�/ٷ��s�MA)�j�l�Ԋ��%��zT�W�J6~Tll ����6�\/zrZ.�Z����-����x�y�7b�M%3�?.0�F��!K?O��S��.��[�R�����,���G�0C�'+���_3w���>�2<��׮[+���˕S
�Qm�y��'��a�Mj	�r���f~o�߹Yl�$���܊f��>_O�g��N���%�2�!����d+W�d%%n���θ�D��Ҧ��O�t�K�Zb��0f�s��8��v� B`���-BXӭ��z�A���;䲊 ������ۥdn�^z/���&m�N�wbX����5ڥ3O��vWD8,�����Gp(6N�3j�b��׶@�f����$������mPD?d"b�'TT�W{�;(���.�'��8��H����Ү{��=��%�>�������4g�G��� jzD�)2�]�г�?
�E��>N/��V�ߨL��8#	ecT�6�rZ�C��s�_�'��=H���~�z^�AsN~���k1�U�Wy�~��Q�U�(iH\�`�����i�2�Â��8�YߜU�fyX�j8Z:������t������v���ό���=�c&���`�G(�+H���J�A:7��7����m �F� "�(�!;Pk���b���p�C��:/�ڏ��6��n��L�˷	w�~i�{��&p4�L���	�P4�p��>�Ԟ�^2����A�){a�Iӯp����NM�
��j��p���HQ�F-�t8�V�wX8p0y�^ZZ��ZE�����J0��N���)M#�,�~q��Ǟ��g�1��w�k:U=�}Y!�r�[s��/�vV����fC����M����}�>����UY�U^�@uBPR�} H��� 7�St�m��._PB��sC�0Xt͇�f|��!�B�GM���3�l^+uς""��57Rߏv|��
�ս��@�Ӡ��/�v�7r�,�a͝-CE�X�" +�qw��6�/9*!1#<i��5�|�}��L�#��g��n},�d$��|�n�i�Et�M���\g�ي��X-�Hϟ^3�')ZU��d�	�<��%��kK�{������Qݘ�s9�;�#�:)�>Эm��4����W�(�㔺�QCy_�;��� J�g8�2Ά��g�gX�}�]����˧F���[��ns,�Y��mt�>y���&�>o����@�Y�p�ȭ>haǵ�U���=�:Y���Y	���uh9���N�?a򦲎�p��|C�C�g|��fQ�Ai�8d^H�`ok�d��>�Lj���i�7!�{Η���Sg'�m��ș0K�#�3�<��C�є�қZ�l[��вR7q��xż���0��PLI�*:֊қ|�gA���鹓��Sp��/2b/����:^`F}%��ا�S���*��QF��\�\���w�"ֻ<�����}u� ����[����K@��J��ظO_������C�֞���Y�xr�U3��%�5)�u&{�Uu���6깫����O�*������V3t(��x��<;�}�o}AE����)$I�h�v���!F�����ĝ�8��k�ɽ�*h&�YYR���ߡRc�CL�x�}O��g�P������j�a5���a�|)�Nx�*<U���9u;C;� �F%��^��C�R
�9�N��Ƨmy�-�Mʶ��;$���0�������HG��5<�u�ˏ͵��sl姕����3���s8ľ�QԽ�̛�3hv,hc��x���N3~8�|�WV���.0xԙJ������+`�]_hQ��6� c��'����ӕ	�p��v�ĥ���wn�b%�/T9ʦ�n�0qB�a�9ʭ8�6��і�����B>i)��]�|�6Ϟ���7�AE/�r������Q����:��`c�h8��V�w�_�B��Mޅ	x����)�&�j��)ۼ]^�4,���M�z�|��*9N�Db�H���!����
P�w����s�}�q�l�R�7ٴ)q��i;�55���u�4��ޑZ?���^v�ř��muT 0	��.��z%{��\�켽�������t�`%Q�}���u��ZQ��ibf���-���M�J�g8Y�Loܔ�V6�,�5��PR^��=��@`�ñ*Z�E��*'{T�M��*~k���|c�e	ȴ��7�S��MT�:2��r��{N.�T����C�����0�W��?���郇�ڷap$%'Y�<�薢�-.˻���w��d�TV}�=d�\s�P� �M&�y�⾤)_���g�
7�$��,��,���O�I~��g�9�WU��N���'��:� Z�aKC�OFhls����6�:'���Ļ�������� �nk6	}I��SG�@�ɸ ��E����3=� �� ^a���<�/�-4��xe���+��P� ��J�emA��o�=�}���X�fl�D)3"�R,Q��������X'Vi���]0�]ѝߐ��=�\;* �dzY���H���}w�'�$��
>
RQ��ch�)Z� �,� &ʉm�]�Edˎ1i��r4�ݘ��ˊm�����U���3�l���~��#Q)��ݐ@����<�X�كQQ_)!�����7Jc�^9�]�|�У��y�!u�d�@����|�N�<��ٟ�ј�@���*��Y���.���܈Z�����T6���Բ�3������Y4s�"(9�$��މ��_Q���7��<u N�mV��1��~_T�0���!��œ���ܯ�&-�>'(�&��m\�Mk��А!�Z>U�y��&��F�2Eq��OMJ��f���s�e�*�\T����ւ�m�rȓ[z����i�5Ó|^��!J^��h��E��l��= ��P=���l7��3���x���>��z���5��0�m�Лٔ������,|�>s"�k&��үy��I������9����7ո{�>>��C�ǯlzY� D2��@��R�q��9���x�u�z����"C�wI�t)L{A��<��@c~9���Vv����2��u_d����y��>�������b?�giWT��$	�-�'9;vu·�瘱�o����p��J��#UN�W�f)5X~P7���>��R���5k�Y4*Hi�<�BE@b���Ձ��3��i��8!�m�2�#5�d?���`���e�q���ԧW��~p�x��t�[���9�]/�e�T��� �%g0���ku%i�Ce��=� ��Q�0�^�� ����N7?T@�����D+�@i�����;?D� ��[��(�a�1	�¢��/��p�����9�u����ҕX�����01(#� !��9������'�O��2�_���ԟv^�2����(Պ�]�h�@u��'r]� �/]_}�y���;���z2�i�O��[����OPi<���7Sx�2m�|j��@y���r�	�jB�ئ���"��O�H&�D�ny2T�/��m��?
���pj|�Nv���\\�D��n���5�r�4�E8L��ih&���+ L���Ƀ�1U�n(�ޥ��X���2@�+�f���G��.�:+A�Cr�͗�`�#�����Ըw���&���ۊ��L]4�i��q����ba��"�K�͡��OT;�K��uʹ�_i��u�#q|c`xI�:�t��6A��gBº�_���q���).(���?�8�m��JK�]s~ݫ{��5UJ=.���/�AI�l	{[�F�up��XoD���q���9��m���]��.K�U���C�	H���N?g�7o1��tC��e��1�!�^��e.c�^��#V�Bq��՛��:0�� �S9�ȴ`�C��mi_��*�/�)@j�����M�<\�8��&}O�n-�h��W���O��[eI��e঱����O��a��O�mz�0N}{�S�M!�{+���,n��ny�0�m�����7��:��u��(�a��gh��?r�$���JhЈ<�M@GF}��JF�a�	�"�zP�8���
��[�t�٘?e�#"�sYڙG�+��jr��Ro�9�I�D�0�R����P�WUq�Pm�ִR�ث���"JKƾ��M�5�)�)�%Ó a) ��� ��1�PFϝ+�*�>�����y�/�vZ�ҚX��Fɧ���Ҁ�U��<��)4a��Ep;�]�m�09ص2��Y�O���s����[��$�r�J�����ɩH#��V�Z�����0ܤo9�vk��(��N�з�V�a;/z����'��i�s��og��견��w��;��#�ǚ0/����&+M ��pH��ы*�
�h훕�Lf,*���c�}��e�ڙ�ά���_���{�<'������L��>CI9��?��|6���^t����,d",�(���o�oq6E��1�c�/tɀ��g	P�:ǔ|��8c��#��� {I��3	�a��|秢�#xu�vC���N��%7���#B�A���`����H(6ϸ2d�|���';l&J\ca��WUq�D�,ZK�����YY�Sr���PR����;hHeUW�2��e�F�r�4v�^�L}
BO�d�Y�|z�>�+!]K+� ��޳|����x"�����8$ϧ)i����H�ֶ.{˄5��5���0�H�m?�����n_���a;�%�Cj~�{s���
��p�ɬ�J�_��m|�o�SO��ol8�~,�WC���z��#䎮W�؀� Z�?���X3�����6�P��ǿ��<��IH��vf҉ϻ�'���?�0�y"9Ͷ9nE%ҪR�[��G@W��:0[���4�cM������5�9����y?Ɓ^�&=r���@�p����ǆ���[������J���`�<�,(O������-���N��œ%b��u�Z}���tl��E����m�Q!�	Q� �	����l����K��VQU�sV����(4�=*E����QV�T��丫�뭐���&�u��v�o��t��	ʮ&[������"���1F�w�3�O�p�#�;�����Φ�JTrE��R��n���O�m:G'6��q��%�m�1d��J�}����M������8�%'�<��bpۗ���.m!t�
�h��x\KQ���wm�JP�u��i�g������`�D�b�ާ:�th˺��7MW�l����!E8�nD˽�H� ��zr�Խ���	£���w�ڛ1F���a��F����������؛oi���$�/_�ۤR�%!p��끧m҅Ҵ���=I����N]�!#�� 7���C��p��;/�|߬Ɂ����F��:�/�+�\p���w��{�hрL��ҒE��m6HU^����ܣ���0�Ѯ0$4��q&v�7��;dc�껧����B�P-(��,H��p�ȳYi��˹\���H���U�;���b�� �b.rI��i��}Z�in���,��w���~�F��f;=�����h�����S�=H|XD����{��0��vHH���/b2ŷ>B�c�Yߗ�t�+�j����x��jUҋ��ϊCg�*������xU���Cp6y���-��J��IP��~�~�B��yk����YTU�|����=t������=�z�f�OS���Y��Y�>�����.&I�2�WX�; �91כwK��X������!Oez�:o�].�`$�`� hoL��ol^t��?:±O�Z��(ciK������g,]�@�nMB�&��������R��ͺ5����M�/���[�{��;r�W��hv�ӎX�4��5���c�7���z7}&�Ǒ�7�ĲM����y��������L7�.(iԔc�'����?���uv��DE&�������i�]�TI�=�U9�_��y����kU6��j�T����BV��O��w7�E7G���su=��!�.��%�����$ʒ��#Rq'�����?$�?�78�=E_��C���B{�� ���*OVtV�dj�
Q��5��n����	��!� /�ykOB�����7���
}�*����$���+����f�>�`�Fp�ۢ�z��D�.5	�Q���3�K$F�ߞ�����z'��麛k�^��ĒnHN�4����6HL����6��'������ս�+���ݼ���p���&�He�A}#��,��r#���t�e;XV5vD������Jt��9��O3�p�y�����>Q/�U�x:N���qJn�XT��
pF ��
<<D^��$DE5�`��o���yY�ޡ�+2�u�hyt�6�r���y�JӍ(v
�X�K��=�f�QVK�7�Nt��~�j���nih�+m�ѓ�S��b�-��Ѓ��
��c���4ߡ�h���%w� ���p��F��+���V�f��j�!�o6�C������CБ����K�����'�Ί�">E+�`���Fc�*���J�&�"��Jo�>�
��w��U�U���~���7	� �����Q?/���_�Ta�r}��	*9�/�5y�i�r�.5�Z��Qy��X>���\i�<@�U@*-<�D#�۴j�J�/��|�n�x�����s[B���Km��p����߻�G��R�T���Pwh��~c���'�Z������3�3u�
J�/*���@���:K���������z̃)����/���˒��r�ͱ�C�u��6�΂�뜂�霎�ÃS�2@k�l��I�ܞ�/�c�a��I��Ǥ�*��]gP��~}�ƣ�t�B9��n#if4��SJ:x��>N���1NU0�8��b�؄�g���I�AH(%Q��z�8H�\���r�-��b�Z���?T|m�����~O �*�<�H��6D��^MӶF�o��� P�s	����ӥ�!�?L�1�S�_���o�q@6-��O�D)�_��I�a�kwa9���.�K��4���a�������D[T�eZ�if���CX��J*F6�9���Y���jR'm�p�u�7Fж�wV�I����[qֿ�AI�����~�V���̈1݉yL�LG-�'
��SaEXS�c�"?�|�yL��A��������j���m�hE׹�^��S ɏ��2ѵ�{O���vK"MN1��Y�Q*�/ڿ�6�Z�}r��H��'�<���0�/ߓ�w��6�IX9��p跉���L/�.�=PPoE�'r��f߂�ٷ�R�=i��k�)�[6^����a�$UU��HJW���B��{-R6-nH�Re6	��8�@�/��uN��V�|=�:Q����Km�pFZ5�Q�\��Ã�y߁�]�7�:�<���{�N社�|��1�c)��*쩨� X��ѳ��i�1�}_�zC��.�u�A�Ӣ������nvu1�托���L�|r(�/S�V��>א�:r>��N��z <!�(=K��s���6k��JRq������"��q^������g�R�iy���^��zD:6�D�=jgܳ9%���_���y`�:�z��� ��9�R�an������Tn���W)BO{�$���Zf7�d(PI܇�|�����������ҝ�a)h���B��3��r��1��/p�	�y{�1��(�/Ȗ'뻷��x�f%Z]ԣ�����v��u EnFI��K`�'V�����H���%�[e�;���\�`%�4_�}�y�s<���2gH�a4��T��S\�4C\L�i�-��'}���=�Bk��i�!�Ÿ���řc*��g��ܿ�����?��0���	����1$�Ȼ������Q���M�� D����+8�ʦ�k�_Z�^Q�K�;�בGA��[N��������˄��uG.�8,� ���`����\�2\1(����E��g��%��"_x�:�%蔙9���rKk[���o�kЪ���$��{r
�~�"`=���l��ٕo!y�?T�=U�T�?�l�o=?"�@��h:������3�*�Ô�#�Y,��$u9��ӛߙM�l�Ǝoz��YG"��.��򋳈�����w�>kf�re@�vc#���@�z蝭O����_����7QTߎN	-���R��-$ߞ�k�S����6�DP>mT�S'�"�_�t�� �lt��Tm˒RroE7��;E�k�P�^��D誢z�\�.X[��x(�1�M�>�ˁM]�.�tU���Q�4�$'
�8&Z���(�����0b�s1n5�nW��rZ�[��0^2�f�w�(j���䯍��+Z���� 搰��"��������/������P����Gz��v��~���ع9�V�j�@���I�#ˌ��#No�,(M�[���/r6��U�pլB��!u�\/1����Xa����95�wa/ğ���:E4&�ݞ�x���G?+^ �=>�)�����?k��% %��z����q%����k��R;�G_����:��.��h�8V[(愓M/� �`ĂE� �!������5�$	�!��.gӫ�Z�ƸV?-
Pҳ9i^�&��	���i@5M����'Ub;�z�P�ͶVI̡K��a�lգϳ�n�%7/V*"�4���t���e�V���f��:�Cb�/�I��*\�]=O������.%ܔ9�����g;��ŤW�Va<]"��_y�c3I��n����D���Lꖣ���-8OزB�uq���T���M��ُ@���1���@��?QE��}[�*�'SrB��;&������Q�O�0�Jg#���I�T�U�%�|��^��ڊ�!��������y>�a L�҇��1kXA�jI���˕�a�/\�Q�a���A�,�1rՂ�g���Ә.`.�o���d�T۱\�J�@�)��Gڹ6��2J]��m��[s����P��>Ir�ƝU�9��0,�s�u�v}n�~��dP[�[�M���F;���W�(�J��*��buV�5����5c2#/'��)cL�|P&�aD�Z6`־`��43o#�U��޾���K9���VZNђn��>�,�2�&��m�*�(}7�}�i_%�'�"ʂ�+���3Y�����*�z:]֥g�MX$W�q�莧�T=y��:�j[�Jc��������o���n��GAu��Cq\_X3e��K��Qy���h�LB_^��M��[}��A�g��F�n�!g�MG)(�N!��ĥ��B�n�H�q�H=s��X^q* �$�.r����5�k���]���+`��? ��~'k�T�ur�{�,"���
E��I�b!��'����[�S]hM�A�j|�.@Hl3#T%�[<���X�"��PR� zt�p�P��Ag�jW�σ��O��ZytH�Ί��C�!�E�w|1�%S�b�ဗU��q��6��R��}ܹ��,�EaO��mFS.u����&�Sۗ������5���ª���G����v�zKui�
���b�5�]���3K�tO�U�xΏY�*��p��u?�����#��AdС��U��)��1#N�=)*�G3�7�=U�X��$9��k{(�,G����d�FD��
��"��;�{�,�[l����e(@����t����Z+�M�gEa�l6@���Q{�&���q��D���7DȄ�Ҵey�M���@`�����>R��Jc%�{z#���*n:	����|Q(@�nLBD�]� ����4�`!�f����^�TMy�3�"�
;c�����dTJS���J^���C�u�z�����cK
ܓ�-�+%(�������.�(��if��'�i&pu
75��@A%t\��0�ӏ��A0X�x(e��9���=���C��9B���I��:ɏ��g�z�)�����W̊�a΋Td���U��I�TnvIm4`"^����I˜D�i'\Ϯ��_����*(�=�f������1��R����Ѓ�|�O��T��[�����-]�_։X��M��NYZ��I1��ۑ���R��Y'=��8��jSI��xx���jc}(�u�B�!6"�����K��6x!�Ơ1A$0�ӫ��_���� ��\�2v�sH�?��~�s���V�u�.Ӂ�q�b�u#J���Ӯ���m��k��'S��s�z�H��D|ڹ>���ˑ�`#�&���"��UZ�VSd�����,J>���,$:z���1�WRR�)�r�U�A3`�'�(N�SPYxy�g�s�.,�l���gх��;-afԻ�H�!e����r��gH�k�&���n�
Z�T)r�:�p�ʪ�G�a-H��Ye���{Cb/��|[-���_�:[�M�N�ג�7�P#X0�
��6$�p������#.��[z��N����T����j#�Y�|њ$>�18���ɯq'&���%`��Tm������7�Zh;Z� ��U���d�������C��� �Ü��173=y��օ�����p�kr*a#X�	D1���ɳ1"�
3P�6��%�����
���h�&���a�fȄy|4�Q� �-��I��A��Ec��"��������\%�}qfEȷo��d�8��%�?5����B�[9W-�r^d_j?{R��=��A&�U�ؗ*��O�W�T�U�v�b���ͧK[btE���H�eIY�B/i-��Ş�+��
	�O[��I�����
��� �?q#֗xH�(�E��'��%��T���WD�)��*�﵁M�U7�n�.����!t�� �9�O�KL����`#Oeִ�p�X�����'�t��rw�|C΂���N΃=��k���2�[���5�ki&��C5B��$aI達�V����������Y��N5�VH�!��6nݐ��~C����=�Kw�&�e���3�5-��>��+m��ؕ�g�m�����b�b1K,kɫW����W�h�B�r5���cd4�������˝\�2��(�>i�G.�@a�̤�|�)�<�jS�+�����Yim]�T�������8�d����K�g�P��� ���e�jԬSc�R0����IR�ˈJ�Ȏ��'���f
	�IbÞ���a�6W�s��%�ځ2Sp��	@�9B!1�a�c�
a��`��o�%.�);v.Tĸ%�����,K-ڠ���j[�l[�Q�7�1񏄅&�*�!��/���</A=v0]Z����;``�8E�����[D�ͻWB�߅Vgl���i��u�iB��p������J�&�%���{YP�1 �j�$�`hu\M�VBĞ��*��c�����566p��&��=+�fL��%O؝w0�\7��Lv���'�J�>gSm�W$ή���AJ������5���.S9�:�5��0}�a�D�t�#1xM8��b��]_(��d4����$W[}��Rn�Gf�*��ٞ�@����2G�$�﫤���_9w!��(O��e��]g�?l�)��:e׵'o�E�az��8i[�9�j]Jq⩧pY�j��{�`"a_��̘;�[��-��o��J����f�$�����-s��t=�1������a�Il��6��^����T�2G��1E�sX_5�&p:E��YwbX��i87�v$Ud����j:����ΦǙ�Q4�5�I����:��� ��1N�A�Y�srQ&\b��e�=�#��xL/�E]����;���7���޹+1�vGO��|�<�"u8��Z!���5I 2��v�^�k�� _M���?��:uL�j�y	"�#
|�0*�]0P��(�]@�;���]�K-a�R�7v�4�It�0?Nqͅ�J�?�5Yߐ/\x�P���I�2bx˄s�|B������3zh���&(�\Q��dߟ�9��L+)˯8��x�u��[���g��♠���U�a�Yo�� %@>#㆜k�WMht�(��$;*��p�Z;Sr'ݴ�b�N�	�q��v!]qJ�aa�z����|�4^�ϱ�,:tp��S����p7�2I��ӭ��n%�La��^&�M�?)�@���.
����q��1�G�w�b��|vA�Z-@�g���|��('�f�������dM�gK_����Zݶ�%�2/G��VAp
0��7?�-<�9���Yn�cx5��"�
V����������XD��qis��$}l�4�K���C�TC�*�غd{O��6���C��_����"}��h��8+�#t襣vji^��T��Ȅ���Wv�����+�@=��p
�O���Ͱ���i���G>9��]�~�̂�}�A�� ������kǾ.5t��-(��*"��֖�|��k��M;'vX��;���_���N����~��]�I�F'�HDYiMn{��@F��(*�a�Kf��� ��n�lE� ���9z��sB�Oy=_]$��`��I��9��C�n�㷖�#�v"/�,PG��@�bZ�6{i�E����'U��#�{e��<�M%�����O8.*��N7N�5�B�Sn���sG쇆��jGM������A�y]a�ky4��~���.
5�N�Y�q�!�~l��YD���!IT*�@��i��)9r����A����k��(�!x�!�F����2mۋ�R��ͻ�Ȭ}���6lG+
dY�B���D� mZF�xt�O�ǋ�`,ܦ�~�y���:
�9��BC��4��f�b�d����7K��0d1-�}٥
� $�e@v\R�J`�NrlMB�;�c�rO_���f�6_<?���q�s��[B��e���e)�K�W�B�UAg��%8���!��*#=�J�-~�l����u-��/J�0�d3y�b;��B�=Ԡht?��L��z��	8����<8�k�Tܯ�*�d��O�L�e�5
\̀�{�<NIB�+uV����϶�-��7��Uڣ�%�X.ƍ���}K:҆H�(*��J���v|�q�7w&��{��FB�� q�?4���	¤Xn��Z���	ؾZ�-��=�.�|:�|*���q����$y�ǃ���G���(�?Շ�LH�7
x�2����ް٥O����$���W{�
�V*%���$�����5��ThbF�X�T*�t-G9ҊT��9�����pꐺ��@�tR�J�Y�g;��z��W�G�E���g������3TK�~��;9�b�;��:ܵ����j��7�+z�[a�]��Azy��Ƀa*�	��,.�^Gr)_l����Oڽ1���J�j���5�O�,A9��'OVn��k�_(0G�`�@q�xȡ��a��q��#\�عA?��_a:���[;�]Sٞ4w�����'P��;v���6��S=0f[J�����1�T>l�Rc)�S�,n��Ͼ[���{݁���� n\��K�D�}(e��1KM��KC!3�,6*ʔCۨ���~�ү���NfR���&D�U�P=mؙ�K����*
�*��Ӟ`�Y,7�#i Y�s1˿[�D	�8^�`��U�V���'�yg+�5DI7�=bR>�a���ڠu(�>=�$&i���9�*8A�,�|� 7t�'�o,��fl1���#���c�]��E��m�*rlYt��砅�����u�^�����uH�E���"W��27�KD�<��v�RzPȤP�!H�It��#��]/[�Q�,L(S��B�[EА��u�z@Q��;Pm�0�_f��1�!¸�ΔeԅY�ߙj0@8�պ��e,��G�o7�t@{��_t�8����s{
A[U4��ע�z)�Fa��p����a��8�7m��q.@}4��t`�t! i1|m� e�q&̗PLի�ˋ]�.�q�=��H54f�QP%���(�E2�J)�Z���C4[b#Gt��C�E7Z%V� �Ͻj�k�QaS�91<����\�&��U�"�CM�}"�{�L�R�/�G�Вq��$E0P�v��Ҿ�a؈5���R!��a�Ff����bB?Rڹ����Ah"�OV�M.=�}f!����*v�H"Q,���G�B7����H�p9����^���Ǜ�, wP�C���@iȠ��n�:˿��29^��k�<<IS�O���^��1�Jޟ���iBmx��Njw;:�����V�^�![�Ī�"��`/�re��P?Pd� x���8�8�N�_�ں*gs��Wh�|�z�+�����4bjp�s�[���8��?	;э�b�ǩΖ�q�Y܀f��V�����!$���+x¤4q���P�x��3g� Uc˟����/�e�ndM��C���`o��C�[�A[�),^j��hZ�}�>���h�0�쥽Ӱ Ǚ��[-T� �π����*[i��e ټ���I��;�z�0�:�*2��ר��@K��g�||��G�8�U>qxɚ���pQ���_ΙS[U wZ	�l�6����O��\�zd�o�DL�#�GT���&���9�%2�"�)P;��؊=�wbRJ���#�\'����9�9���E������9�T24�s�����êD�{�i�.�vTs("�z��Ct���H b!�[�{9~-����L_��=]˚��F�"p������o)���ܑ"�z' �'o|mi�)6/K�q��/��&�q�0gԁB���.�O�7Y8xr�+���v������Ҝd:,:�/?AC��d���x���9*Q����lo���#)����ʱ� :�Kqy���cw��}Ӄ�zY�\�ꮫ��mq�)�64��bP7�
%6�P�Ē�/S�P�{W�*��}���K����:�����,�<}E)��n,v"���hՊ9�n:�0��;t���n�Q��v$,�Ǥ훞���S��e������H+�T��?_"���DN҈H�`��O���j�BӎSi�L�I~}B>�ZM1@d�>D8���,X �}IyH�&�X�?��Q��l�8:/B�Z?4���o��3Ʋ�7�7.��p�䅃����󅚲���J�.���լ��ǹEZ"�h��FB��Jռ.u#P�U����G�Ϧ�t��ؗ<C�mV�j�~f�V#����u��LW7�iY+P9�w��B����(!bd��~�o�rv�A�+x��%�ѕD�gf�S����p2���Yg�ǆ2���r�m��04p_� �a��1CTՇ������F�����6,�J0�kOL��'0gיg���YG�k���h�5D�5�Jb�T�4���;�7�gj�@#�ͦ�'������ r��{�bF.��>F�Ѻ)Gf�{��N?��9�Y���ԞJo�\�9��Y�Vr���V�N�P�k����=�Uܠ���w	����'��������`/�������L�Q���q0}kn���Ǘ�k���������I36��$&u�2��a�m�_�͝D�a"*L���$�ˌl�C�X1w����}e�w�eL�OeSJ�@�H�x ,�qV�4ҥ�9X����в?F��O:�3��a��.D[�U���)�f&�i�V	��d|Z@��H$���β>�qa�ATT��Њ�\"����swF^�}q+����&W�E���?�]��`{
��wN�L@��,k�Z!^X�$�K��$��y��3m'(?�&B�]�n�V��ĕ�z��L虃��D]@5.�w'��� �޶�	��^e�¥D\4�o?������?��e?��_�XVߗ٧�%��VSX^�L��]=�O@���,n��j��t'r��H�(Vo�ƐW���;�E�e�Ȁ���/�c��������}�;Fn�rP�y�[��T��q�w<�
6@ܴvDy7����*������ȁ�UI��/r|rC�䴛}R�8Ι&/��!2���A�Ĝ��XZ�|�"��⥨
��IX��D�}��yP��V�{�>�0�9���w0�����r W^����lN�+X��V�=k�O8����i����ǀ��Ĕ���\�Jډy�dEhtI��v4tġ�X�������oM3�ŋ�4)"�y֖W���:�������5P+l]���ׯw����F1.*�d2��̬"�kM ����������y�`Q���%��9c���Ʃ" ���7 �Z�k6tf"�������ɉ�5�Z�.$���%a,v0���J��v�~ z���V�h��=�f���ݤ��{����	��=������LJՔ�ˁ�w#�?�����V\n��u��!G�p,�n����>�@�@�#�g2eC&7�ב�B�����M���k��e�ۂ`yGjh��Z'R��y��PH$l<1~_y�쏂��ʟ�^�R���+�e9b�%K��![C�P�@F%�����Ca~���A���KJ
��!��0)Y����=��TR)hJ�0ʇ��j:��O�K��r[���/Y��b�Q�B������j�6�������} l�f�+{}�In1��v �p#�+4�:*aP���&=��N���n�ÓOB+7F�=�h�=�L�o���o���pu8BG���I),�:�O������h�tM�×4��H��K�GJ��R��vH}@�8?��Z,/\�xlgd�_�?b��5~�����,K�1.Dw���#R͠�����
�dU츦�Ӳ�^��1�	��ֆ��(Ȟ�%�0�J~~��ܹ�~RA�a���{��$ $3CdlW�{PNF=b��_��d�by7�`��7� �FI�^�H|�I�g���ou��-�I�0�iyU7�j�U#�����R�������9w����|S-��=�3��p_�)�o|�� ΞuLs�8L@�)��]a�-p��1d�`L�yL�o@*��ȶU���Z���˺��\���P"���ObևN���3KKo4&�L\Ϭ=�S	��Yc�?���w#3W�3c�v�eЫ �> �>�A�9]5;��cdK��}����0p�o�Qx7x�MS�] '�iS���s� L?|�Op�n���5v�(�Ǆ_I<����80͏�5��ҥ'��p3s����O������(�T�>i��jhƙ�'(w���'+�j; ��E�<���H����eWa�dLy�5�I(��(g�إ+�A��vߜZܠ/m(7i�l�����[EH����Q�ݐ�:[���U�YQ*�r2�D	�Jl�l�&���t�j�"C�+'1�����l8�$�`�����KP`;7A8�QΧ �1G^��y��Q�wA��`�Q%�$�h�ס���6# ������r'VAuG��\sT�=K�Kd`�KX�Ų�I�o��(%��,d\���TUͭ�E��'�����J��x��D��T�\D�(�?O�|�/j2�x̯��ڐrpb	A�5*X��7S����~�7Å:��"K%:�W�������?#�������l�
YltO��0'V���~�Z�e[D&�Z�|�qɍ`��6��X���]�i�K� �l.8�����y��A��� ��&����~5��.�����7��Q��s �?�y�Q�a�Ǳ|��r�;]�F_�����%� ��|N1�s��A-{@��^��������&�r���>�2c���=-�c����rM#�/���Z���a�\2�X>�ivi�ؔ�e��F�
�zќ�.��J����I�i(��877p�3	%]? �NA/�;��ޒ4�W�+-Q��:gy��+ [	+]Sm������='x����kT�o�۽�*��������/C��5C�L��A���+gF'�3ƥ�NH#��Q~j�_�\6���Aw����]���:�����	,��� i���x�i��灸������e��Ї��F��]k;�w�n[8B�`���R��[/>#���#�s3�֍Y���w���V/�7E	޻����d$9����@*M�
E$A!�ѿ�x�'�o�oI٤ִ������ȫ�o6�ղ���}�W��:Q�9�`�R��>Ծ��U��j�vvY'7`I]N;��ʭO]>����F��6�F0'&F�:1GOr$@��C�h�%3/��'�M��{f�Z���9gps�Po��c��;Vbm����ݽ=�dx�M[��W��)��酻�+.X�������:��z���2M|0���͹�(��w��T������u��q��VZ�_��t��8�M*�� /��\�'�3���E�I�(I1#��R�c���*�O쟬��,��e�ޣ]��|	y W���n�3A\'�1��5�L���/e�y�ŏ���w�X�0W���X�/���Ga�<�G���ߚ�s{����<���A;7�q�L��-q=�ةh(�;El����xC�<2cC���d�GT*��\w5��q���h���B׍�;3�@��H��Z�a�Z�;�H����|ۆ�D��
@ٛT�ʠ����M7]������ca[q�VM�P�l`�4�I���&�$�9(!�8�޽�b�u7mد8M�(������4���Q���7�\�z���cD~�s��.���L���/fi�la�� �|�%�~swUG��G���o�XhΆ���0:��N�KD�쇨i?�{�Q�?q�a���6��d@��n���%�T�{M�4bd�Z�=Jy�+4:�?k�o���B,�d8DfZ_hF��Y����k�@���F ��}�]E��j�g��,���Bh��B�خ=�
i���N��� ��P<�`�L��q��E�ЈB)=c
��W
O#ڢ״QA	XYɾ:W���@�ĉ^�=A/W���.����E]�M(�Tǎ��3v�!#z�6.w���O&Oi�?��=;&�c��8H�Yb7�W=*��S�y�V��2IZŠ� �>��ͮf�ev�br�����{GiZ�{P(�0�-o�e�8vL&�B䤖�dh��E;D���M�.&��"�l;ViL�v�1!�Gi�(\f��;Ɨ��<==N�B�E%[���a���&$���i6���6s)�D�����\09+�(�CS�uo��Q�;��=Α,�`?/9jFq��W �1nִk[���Vh�Kx?�DӪ3x�0J��:v�!�xB0F���1w5�;VM�;xy����#��~,�m�/�\��Ek3���Q>B�б�ת7mi�7�``.���p��2�>Dr��; ��W�Dah��	��d���Q���Cù�hu��p�]�C�����B��)���D�,�H������N��J��ś���w��O�uX�8��X��@R51r�`�WJ �`(���'�Rs1���QL���.}w��4X	Y-��b�~���!��}n��ɖZZm�6��q%��Eno�� Ǳ�v��\5��B���K��k�i����9Pi¥inHr� i�E�F���q��5�$��yK�<O�A�&r� �	҄��{�^�~gm?�yQ�ޚ��2�C�v���O0N6��~���jH�SD;����K�!=��^A�&��	�)��@��}8�
�68R��ߒ��x�?����l�!��m���A���A��G0����EX��)��C���|3P���ݳ@����:*���=� =���w���{Ҵ��L�M�z�UC���+���ƩF�p�a��B"�b�ذ���B,}Zڃ��=������41�9|R:���32�4I&Z'x��
�El��R�G�pB�i4drҗ#�����2 ;j�OPgFl��f�y�B>T)=��K�;�u��~Z1T�Rk���%���k�G���<��>N7�����.�{�:�G�UIy�E��VU*ZG݊b��yfA`K����7�jKҟ��jL3^F��-t�%y���� �2E-����m䆣� �R1�_t�]�Vel$���#��[ߴ��4;H���D����Ս�T���u�G<:.({=h��? �I���g.�D�j.�z�Y){o�i���{���p�2R��lXi�|�i�PVܶ?D�
�`����n�-}��-|P�0�x�J*z�Zq>�*yW�=�T��#�z0jk�j�ʥm��� C,��p^�wna�h|1�t�����1p�s3ظ<q��P8�r���r�RD����{ޔY�ܴ�D�m�m�Ҷ�[#��}����Y��
�Źfh�6�g���Ya��l/�ju��ǫZF5�|�1넛�*'���֍V՚d��Kv f���nLR�{j/�i��wJ;���N������0�^W�%d��·+8D�x
_�1�V�OYk�˹�ExZ�Z�-�KȦ"P{�V��� x�!���p#>��f{�%s(>���BD�M�#��B�~�� �v�sFV�'(������	��'�i�{�Oڍ>oƕ.�z��	�!�q�XE!t�v_e��._TD��b��F��tO�Ha���d��;$��N�ӣ�vܿ����XC}�O.�h�ߡ�I 4��YEʀWTj�����4ﾶA3h�<�������Q��E�s�wW+���ϯr�q�g��X��G`�|^�@;��^���Rn�	&{�Eo�_��WYkq���֬5���� ���E��3J�E��}
�Q��(�F�׍GG�Us����@1���o!b,��8�s��K�?1q
/��rMI;*�k��b�!o����R>�f*��6#ˋ�v߳�xͩL����9=�3�d[#�5��c�!�#��Ey�W�'����U�A<���f�~���pzCU<t�,d.�2n#��FW�5Dd�b�h�N��T���9�fJ�Z��O$"0�5�ewjapG��"��D��`_�l_S��|W7���)���Sp��u�*�m��tN�P��
Q��-�E�o��1~������}��ʔ�{�V�ĕSF��I�=�dS���ԼA�yj���#��9�1��c��8�k�}����j8!���0�㤝_T��F}�����w	��M�YeOYeA�XO
$i�I���~��`�1�c����&�n՟��������s��
�P.�~~�C8p����)����F�b��v��4�2�{9t���Q/J<4.�Q-�X۝��c�t�"�����+ؚY�B�)��kPLf�}����`���Op'\��O9���hL��s�k ��� ƃ��$��{W�q��y97Y���1J�&?_r��H�=:A3�I�`�c�5n�b�0�q�P��)����(#3����R����o��~M�Ȟ��z�Z��%���"=P��H,~�sb�i3�����<v�=��6�i�%<�/[m-VƝ��t@�[�zv���;��;,T��'�3#�7���u9��۱11�?k�U��)�z��R���W�`JԺ�@H��a���u��~�8��ܬvG0{��N]�@۹p"�;��4��][1q9�nx�=����ZЦ��೩��4#3�-ӏ������y(t�װ��X_`|��G@2%�-��Q������F��+�Z�ؐ@N��s�::��M��{���\mz�K���B��[j��(�Fz��}Hd�£=',.�?��)�Wzf���-i�X=jo�H�'������\�Xߪ3�9B��!��G'���gv��'wO�B �����k�A��}B]�n��)Ϟw�p��A_E�!�~2�Qe@o�r"F��.�E�MW�g�{>�BMEk�f�fL33�L����4�+1����Y#7�G���'��>�B:~N��W�S���	�H1��n-��$�5�^�n�g�2z}�2h#x\
��'O��8 u%~�ai�����G�;|�]$����{��6�3��3L�0��D��09�2�������Y-�,����=C�wΤf)�/�G�YQ���5K&�n�VV�0����,W������Lw�a|%*��h��y�Z��Q�
�����&�P`�f���ə[O2��S�#�8�	&�������v���{zo�b�A�5�3���b�G�ꎳ�"�	E;�6 '����d��?�^g&6��	�Z��0��@��@�|��̛ �0�wG 
݅ �����ݺ��)t�����lE�� �R�R���H��>�?8L�o9 _�3�F���H� xS��L�q\6��ψ_��u��ľ�2k���~oA����4IA`'"�7��?�)Uŕ�r�����z���!�'�-���'�EG�[腗���J�2(\VF�~Ͻ�/��vT@�+�9]�r=�f&��z�'� 	"2j�Q�ǟ;����;�fu6(8L$	�T�T����(��??��Xk��Oq/��:{�Ch�?��au�����`@��T
���u|Oz/��Ǒ�I���C���ChM�	��J�����'��`�Z�ꇗ�yr��4��(ΐ��l%��Bx���\�'j�&q�M2��jU��m&a]��ئ��󆰢ER�<�� ��P>M� ?��&f
���e�`'�-�:èp����-�g�*�2H���7i�0������hx�db����;�9��ߖ$�̢]�D!�����	��@�(�����T3@Z�	S�I��JO���Sb� ��(5�e�	
K>�,����[�`iO�l{�ܼp'��~΄�j�8o6Z�N0��V*��AC=ܪ��O�~^�(8q�6����p�/tF��lgo�|���"���}VWќ���z^�_z�G���i��s'��̞�L��P)e3�H�pLL��94$P�|�o����C�Ʌ��h)+̄��̬��ap~ZZ>�V�����K%Z;��o�C�{�>�2R=2�̵����[d���7QxŰ�"���'��~�����	$(�ָ� �������o3ϓi����,w�9\[�u&Fx����2z�����1�3S6��* �Sz�=]�-��-�{w%��^a6�^����5v\j �:�Ǜ�K2�B�@O
^L��Z��й[�R�D0�\��=�Te)f1J��p��*�y����e'�rLl�p*�_�\�HI.* ���W�vL��b�!������B��ro��I%���E4��� �a��	�8�����S���}T.^���$�T��׭��z����_�ݑ��³~O�� ���;��4�6m��)���%Rq0�x��Mp���c�X�d�Kh`�)Bڱ�\,Yh.axS���
z��C���	�rn�| �J���*m�_T�$;��$�Y���[yem� ����ݻ&ܦh�~ë'y����;��B�>�7�Gg��Vf�g�ɱ��vQ��П���QL���\�؀<�m�C��4���^����t��t�6�<sˍE�G�!Z�,s���N�7֨�V+·�A�2?���@Y�E��;��mgn rc�X�`Qd�$s�4��Їܛo����D��5�&a�_xZf��!2 x\���o*�3�I�g��
fS>z�(
��_|�|(��ʿ_S��[I>�����y!���n׊����PH�-Vob�Z7K`����\�7����8��F%��L!N��*��E�3�q���M*��\`ef��h��ܶ%n|,�N�M��b��}W�%T��g���6�ϡ,��U�7�s9~�����n��rp��Q4W��3m>Մ8�[�_:�!)�:�b����~o&��Ug��f�Ǳ�I֤ٜ{4@���r��1.�s�ЄJ��,���,��ނ���X��u�����O�*��mK�ꊍ`�4%�!NNt9���A4S�m�)��͜*I�m4�'��N��4�9Kط�4�Vg��p����^�S��uk���O�ƏP���r���nZ����`�
r�L��f�c�!����
�uq�7P3	6xm����=yp�/����C
#��,�BӨ�	�p��y�S&�E,@d�nH��b��hJ��v�+�5�"�l��lAӍ�1���zm��-�󒑙M2��˭;��bЇ"���-(P8M�uw�/�| �;E�U��{��	Ѻ�,�jh�$G'x������n�g�ي�i1��Kڦ^��k'˼4��"_WZ�vp�B����7m?J�1/Өi��o���L���.8����pFب^�d��ԃ;O�$כI��\�޼&gE�uN�����E-����*���I��c~�O)��ԃ�E��j�8Y�ӧ p
J�K�e+��sbL�};����9O�����<x���肇uY�3)9�r��3��UK�V��c'��h�vy^+���+��R���B���j���mG���E�NEZǶ�e?�0:+����UDٌ�|}" cmX]��%�!ْ��:�h̼ëB	M_�k� ��N��5� $�92ѕ5ZLpX�>ߐ������\ycx�)6/�O�xR]���Z����n��(�N~�����+L� �B�V�1ۧ�Ϛ�@ol��J�Y��E�6a��:N�+�oC�r�~��6����QT7GyJ���`�$���߹{�^v���W�ѵ
�V��Z8���|��'�v$p�w�S�����T+��Г_��Φ�G��NP��,ĸ�O䦿ގ����`�^��6�4�S_%'��@pWO0r~���E�1)���ˤo��$o>�v�WU���4���;�O��fdj��(���ml�E]��X�3�`�i��-��ɣ�����rN�=K��q�X۲�R��,��|V� 6�^)�o27c��x�S/#�*�B\V"kٸo	bKh�����k�n1���v(��4���D��Zdһ��n����Z�?�QP0Zo(��
�u�䧏�w䮿(H��bL��d�w�����J��h4a��*�k�A�N���	�B0W}T�Sɠa%�{��r6V�!����������sBg�����䬗t��F�dhP���̗ϬkR�h�hf���n�Q�a�n�=a���N�.��@
=:�Pj���5w��&>nS�_*0���&v�b�Uc[6���`�#�aZ�銔�b��ɘe�Q�?�n�Y3���i�E+�E6��p�����b��r⩬�N��\���v��7�H����c�;��3Q@�'g%5���
�)��l���ϧ����S��|�T+>��(���v�4��1�
��ğcn���Kx_�E�(�H�fmS�(�:}}1���|��wy*�ٷ}f�ݢ�@�=�s-�lsL6d��wp�N]��0��S��ؤla��A[�� ��:O�,Ik�Z����z�ŉ׮d���"�]o���<N	G�A�Hv5��Z�mo���
Q]�"{WY\�3"��v�定�=
��\[�
���R&�I�c�:�
��������Q�D6�ϧ`�k�����N������[N���[Y�"��E*�����k���+Y�8ة�D�k�m��UU'M���U�p��_.�fzO1���G�O~�M(Ͱ���&��sNTL�aשׂ�X;.z�!6j�����H�P�{�"��	�R�=��	��܋ib��������%'�v�9� �HL|e��B@v�X+ĝ�*ĉG	�E-6GleTK��<E��N��Vg��Ȳ���uvs�㮱�a�%y<g�O�
-BU�ǲ�"Qu
��!�wB�;p�`ǐ�EN�`�.��/(Ë�����D�ݘ~�|3
��,��K�� z�8)⸡~�	����O�
-�j�l��V���@a�k�a�;�<K���h�6���;�"���M^��T���c��={�9� e9��3��M��Wb��Cث�I4��M�`-�j�wF��R6Jm4���{�ͷR!�>��q�[#�����4l9�~�IϏ{��Ζr��$�<���
	�/=�r������l���)��m>�\v~x��C�+ΆFwÇ7��(i�I�wnr!QbU-�q��&�����xEpCoJ��0�|�S�/ @;���	�σ�F��ۅ�QHæG���xnmZ�/�d	I�/F��I,0�js�;G+a��vŚ]��Ǣ$K�Y��fƃ��9�����O�A`v���"�̜+�J�	1�w
Jt���*x	���B�3�ΧC�
q��_����UO�}d5yz&�����ކ�N
#��k�p����U|���	P�&��-iW-|d�����	ue#d�����?�c�g�'ޗ�#��~)�l����唟8ʌ.��$'77B7+~/m|��.uS�g��@�軅G��I+�A�5����	_��dj��T����Xk�#��_{�6Ι^�ڗZ1�]P�W8�Y�w�z9z��� t}��U����.�*+�IO	��a��d�p��>�.��S��/����ތY�^�Cܐ��c��c�O7���zj��k�qM���3����MT�PŮ�9H=��^O�@��*]^8&�#�a�Tc�()��AJ�vn��N��O�HPF���7�Ȼ�qBg�f-Ź��2K��pi,��� ����:DX�i2���(-z8tT�J��Pl}�PZ���>�C�@�HJ
V5��5(W��`���q^����$��ۢ��˽Qh�{�L��5�����7̏y��3b�SN�_R����q�[�����S��0!b猐r����wg��C l�Eͤu0@?�U���i�hUv���w&���i`�ܺX�:]fו�0<���9|�����]:��G�G?ؾ(s��B��W�\�7y�&ww.}=ӌs�)�@�K���R��Xb�e�_�21Bj.�g����o�7�88d^���U�lA��v��Hz�x�:��b3+���̭Ih��`S�ډh���s-J� �vQ&���h�.>�1�#��́�DG�|��w�W_�@�&F_y;��7�CD��S�c��_|�+@qt7���pW��W9S�؝�/���5��A��	]=ܨv�D��p�T�A�p������b�t�1`D�����5��N�\���H}�*�dQ�&�%gF��~��l ��;V��ir��T�AjS��J-�#�5�VB�w�ǣo���7o�E�ǅ,�#���d+����,�r����'��>�[k,���D�_��`�K�����L��M2Qs,><��:'Ky�����0ֽy��$��g��?�n��:N.]省�N�Q+�>��+Z޲�HQJ���  ���1������9��n�-�6�i�ksC���KCJn�j!��?�7wU���ކ��8��_)�RtϏ6�����N��7�[|�֙���Q�')�9�t��*����ݼ��.b&k5�LkF�߇����thb�<Z��Pb�"f�?���=Ê����O��Q�L��C��1��J7��-�^z�9C+�{��w� ��)~�÷�'xlivD�5�ґ˕'�lF��Rc�2m�G8��k��T�{��@��1͹��R�ќe�ޑr��e�н��m�Ԉ�'�g��e)J�nN-Z�?!�0V�f�UJ������LѢ�iC�sN*?�g\��&U߱M�a�F�Yd{�5d�Urau [�J�h��	�p1�w�ij���R�{1��}j�橦̊	\��n��k7/Q��1���Y�P\@p��v��Z�gy��+<t�a=.r��#׼�0�a8(�'��ٝ�C�9O���%��|���c�pjH�p��C�Q!��~��r��6���P*�e)�3��A�c�������l0�a��΄�8��%ZO��o�����jP�e÷��ĥ�Z[��g�T��u�h8<1	n�4^�|0e��m��BS���L��5�QAѩ&m`���U���/f�'�^#B���VJ����'ĩ����E7VB��������L�Q���#�����*Y]N��ًf�W'U�r�,j+F�� �Ȱ�w}ٞ��M��\��5�`����Bbg]�����4�U���J�h *�^ �e���%z�ƪvc��:f�>-̛��f$�(��w%�:�	��RB�H^@��u�A��vv�9c ww`me9��6@m�T �}"���e��!"������5��K��e_�b�UR�� ��J�ƛ1��y�u5���.!�٭x�~���;u�ri�'�x��$�)�[Uʷ_[~����*�3l*��
�^�n^q���	��V[2ih��XK0p-^6+`�)�j��H�����k�m�~�tK��^<�t���>,~�7������Y[���d�ك�6����5ճ��T��ա���USI�u;yS���(c9jA�֨�.wVr�=��{�J�@�U��ت<�g����Agv��1(�o���2�E��hr�����Q�CLO��ڌ�A.���L���c8n Q� ��TZ��'��չ��(�K��JM�l(.u�՝��O>X��zJ�
k|�ENp%ҦfA��
�ȇ�2���%�<�'�_������"��ԏ�d�j-��9�E��U������޸ٯN���#$RP|�$\��8vhyty%h��=ȭ��n�R�^a�X0������=���p]j�&�)�<���T7~b4��P)��،fz*����إ30$�覔h9K�?t����o�����YaB�6ʠ"���S;B%�0X�u���B0N�`%j�b�uI¯���@��[<){ឭH����g��~@J�(��neC1s�(�ğy�6���Q�M���K{}R�Wl@}��6������꺇�����\�d��*N����U3NG��s�W��Y���gXu$�K�y�lDj�[����RĲ��MZ�h~�L@<Q��`B�zEj�k��h��c^T��at�!������?��x#z_�0 wt���˕�F����}W�x9�����k���qk��o1��aoߒm
��ip#ǧ��RL[kn�Ƭ�����l�X�?��m������<��v�s^g#or��|ѻ]$���J��lO��G	��y����"�{�1/�u���jg~���t��|��"j/ȨL�AM����*���V���u������;��]Q���(��;4�.4�LIV��X.����Wބ�xQ�Z�ܩZv��c����{ʣ	��35��^��E��i?��z�@j�:����K/���|���$y��߁��7����(�^]���e�}���|�KnJs���&`{��V��/�������ˣ!�7wh�0��-�	���m_���؊���Y*��)����EkR ��L&���ڽ&K�%\�	����v$=&N�i� 0�&��Ά�+���b*�K�X�lU>b��)l��m1�[t@9/��ܳ9!�jO�[%�4����l8ew _���[Z$�.)��t��#��(��Te��c���N�GI!m�@�..��I�)fP��Ve����izte�`m���Y9$��P�����R�V�t"��R�142��*p�����ɻe1�vf����e���ZXS�<�s�S�zpU���i��]����������t�jO�x��b�-�R����uR��!Bt���7@W�v?q0���(��=�2��9��n����ې��͝����KFq%gjǛ��ZC�F8 ��N4-�^?���n�����{��5k�^�_&+5أ��I$jˇ[��c�**6H0�ת�-���Yx��Kb�L�o# 䤁]��0�X����WV���S�?"	�`"w~�x�.1�K8�H��@���x{a�� �-�
���;G ��܉g"�U�Az� ��]3�X��9�W���qc�6�����Z��MN����ABԕ.��c<�i�!K���V�f���Y93P�БCVC��^��!�ޱO�p>L�2z2Z*�e�(�')�@
p�M6.v���{;@Sff��5�F����n�Ȩ[�+����5pf�??��ϴ�?�۟�2�O��,��pҢ��6nqy����>��G�+�͆;N~��{,�2c����?7�y��(&Za/��Y���@e}F�=1�� ��Oh��3�s��§�
t�9����XOd�ղD,�rE��G��^�'>v�6Xd�H�z��M-�o�]*u�-��c�5^Čv bT���Ӻ���txRl�Nb'�9�~�#�I��R�F]������ld�x�A0�a���(�+Y����؜�\ �=����h�e�0��ت��4`��3���UB\�q���h9��g����D{R�qH�!��;���u	ޥhC����	Ψ��'�u��rq�u&1�;�i�D���^�e�/@�A��������u�B4/��I��x�{����b6�����^�""5H���^���d�קu�� �$��Y,7�v`ao�7�G��K8Q�"�tN�h/b:�J�)�&�d�w=I��t/��=�w�)���!Ĥ��I��7�V��T���o�s^D��Znw͍n�Bq+���`�fH6ܵ�U���@�ٔ%��'Y'���|��O���Y#��1�H�f���'Ȧ���%c�#�o��vF��`�PK';c`ę���E1?ln���VM䂼� f�����|V�ʷ��5���p����xԅ��;�y����.���B�"�2����r�)mt[����9$<�=*"��
��zz���	���i
~0�_u�0. �oٸ���kp�V������p��� 6���r+|f�~u}6N���X!>Y�rM��$e �\bqi�RS����-���)��R�R9�u�S�[�F`��s�ZH.'ߔ����b{�c|d������8�)g-۟�TO�
+�R�j��aP,%7����M��Sh@�_��xA��r�rN�`�u���ņ�%�187���X�mV�4� ձcr"n,�7M�������#�p�à�
\��n(����§�&K"~S�+
m�L=z��}b���$�����kEj�v]���q��f=��� OW������A��b�V��o��3�F�����l�=�״)�H!&}sd�[�s��ѫ>v�����w19��~
�����WߣY��d���(,���{=�>��Sf^R渗RF��$@�Q=�F�
�`5�v�"�Ȑg�W���-�I����O-� n����ı�5�q�y�k��]
���>���ژa5W����EBo��{*�V�G0��5B��Z�-i�!W�5��g�j�`��-(o�7�LӸW�����r���v�d7�z�߻ue�M#�w9��N�^���"�gw8)��ڛ��2����Y�[��C���j�$0˦5Sa=�m��/�uJV����2��K�Y%<��kx`��3�uZ0Y$��n�>��V<��	��Z󥳑�9��ߝ��l����颱���̎�؉O�I��48��j�����]���!m�]���R�6<��f�}���q�=S�6��A�,�q�(c� JC=2�m����`굲	�ۚ=�.h9�؁�.�G8�P`���&|��"�֌�.�*w�|��|+=1v��.�~-X|�{0kɩ���A`C������,6��f��B�n7ҟ�9��Dn������]�^&�d��;m�@�#P4N������r�!D��!9�r�T�(F�8C�{�l@��v�H⧻�������s��2��A�4v�9 ��fɂ���
�ؖ_�d��^��_7	����((4�p~|��4��/�rD��۾�%���(D�Qo�a�#��3
AXy���ϕ���r^>,ހ3��X�����0A��A���r�S�c6�
v~�O�XMw�z�	��n����vՏ�a�?V��`���W�u�֞��]�)\ Cz���՚0����s)(��D��FA�FOrP�I�3��ٵd-�X�DU��d�<V��#�T�_�nN�:�Q3c{�O��w��ς�[��i8~K�CBD�}B!`}Syd����B��Aa �s\�{fZs����m��!��%�i�ҭ���o�A�L.�5�]� V�V�>!>C6���fؖ٬P�R�&��r��DD� ד�����9C�E�UX��z�	�`��5�ca����f)t@������:�7�KJ����������&�/a`x!�]�1��?��������7���N�7�[P�r�}�&���Q�n4�����)�0Hv0�o���t���L��܇V7�D�4H���qr	���	:3Q6\���y����3�f��Gޝ�G�z�/<��X�M�hUL�Th�K��ƚ��ENg���b���
Pr��MFfw'��L�����w_ؐ�5�� ��-SC�A��$oȐ�&t5�$F�(�����j�������cAq[P��@"O���b��K��r�7���9�w&�N�d��Sz�b����[�$DO�ua3*!��|�?�K(jתy������&|7n]��$Bmhx��	�&:Utx���8(��;��9��|�aO�+���|}x�e��3�X�ܰ�J�p�b�r���q$M���]�y#�q3��	(7K&���Ȩ'ݸn�c���
^4���� Ŷ�5�~h{��ZQ�39#��-�T�+���������_|�Va1fE12�I�pcA�n�O�4�d��A�9T���k�s 6Y�.�n�Q�l�v�)ͬ�!i[�����^� �K��A����ۚ��=6�]�&p�������F@�8��.���cC�k�~�7��ie�x�,�~����[�e_��qe�D0�'F�<��T��Jg ���~���Fpe����z����	-^7�v+I�d!L=��ذb#���4�i�Ƒ��!�)� e�����Q{�B}�N۹�o���V~$����n��9��v���c��C��#��*r�qt|F�| ���_�Q��/��v��+�A�s�Z 2�S�8yX�}$K7���zW���>c5��J�)�q_-RL��P�L�M�K��CnL��Uϔ��B�{M4'��TO�����e|�K�O����z*�B�Z�#1�
[N�.�pO�n�}�-��}�#�~��$��Y*��%���K�ٞ�.aN�fHX��+Z