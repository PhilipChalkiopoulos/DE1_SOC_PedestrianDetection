��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b�������Pp�dN� �T
��l�S���h��UC;#u�+F�p^<�F�ƫ�����V��]{��滀h�&e�ycz�C��/T������1v��S���	=���K���+*E���8��b���I�J&��0o�6�45�e�����<�A+we�����r �S�gE�T�C�b���5lD�����A���}�]�;�_��rJ������UB��5����"M�d
ϠU���C����9��ϼ�-U�٭cL�֚�X�m���wW��N�,�����{8�V�5`C�I�>vdy8� ���e��������C�%�~E>&˰d3%'רՀ{��}�¦��4��r�=�"��_{�"xt2���]�>���N��yF�h ������;����{|�:�G��&D���t��!�z���E��/ٙ�&N��m!"��*5^���3����,Q6s.��qAي'���J��FI{9ٗf��IBL�وZ�����z#�k��[l���=�G u���`y9n��4���?6f�ń&8����t�*����!��~L���?'��Z�j���U��� 
=�����lMP�
)lX���:=wG���VK&��o'KA�מ?}O�m����a�0������Lah�ܘA��e�K�f4�" �3���N/a�Pa�����7��ɐ^Yn�@�FE����G����&� �m4ޝ�����©�.@.��0��m��G��H�=\�e���K��D���m��pF������������ jM�B-�'K���G%�C��ݡiB��_��3�N����).��
���,P6]Se�Ѐ����8��K���������{cئx���C3���ᬄ�+y�ß10j~ (�W٨p���1�FӚ:�!ʄ�S9� �-nq�U�]�	y(�h���LEq�Z�R��ş���_��3����8bC,��m1�_{$<`�Jq;Zx�kw��s����*��F����O��/!&��r�eX$;\5U���y\i���j�)�b��֓M��Vg���H:�æ���P�Y=�]pv_g��O����`_��X�>�3���A!��;H�G�N&;��=T0��N��$iE����&]�����w��(g�GC;�rɴ���]�e� ��[N�����&��0G^l�����G�,:�P�V`/� I�q&,����P�������ȱMR�ocu����'��;�����+8�1=��C}IO}j��+
3\��P w�"}��O%���Ӹli�j��u���U ����pd��J����N�	���!�h8��{e,�l���=��9+&�q�<b��/����
��n:r��%��Qz"Lvl�ķ�~�����w�p��~�<P�ͧmB1f(� �73W��
8x�g���:��Shw�&z�@pJ��/o�����k�i"|g��������߆G��v�O����0��<�}�:~f(�U�n��`/�E|	/����iV���he�h�Z�_�i	��qoa0v���1R�yܧ$�;Xm�_F>z�}� M�Sqo�ݗ}@�#�Aa��=�k:� ��/?ޠ�^O4f�	�N�j�kR��tŘ��$pL�AFZ�V���ҭaL�XR��൓��`k�ëx���+�e#�gT��~k`C_,�AXH�C�q6)�ۉ��F���N��ѽ�|Q{1W�EgͲ{��� #T�)��_�hpa,�֏�jW�k�,צ/��U��, �Ti4�T�g�F��F��dXj�"����_ċ�
��f��N�#g�%�Τ��إq������ H;��%$�$j��]�[��G�l��14b��I�~�.���P�=p�!D(���1:�>7C��$ew=8�c1��h#�����6kS�H�!4��?�����ط�s�A?���@��!��kY��_Y�K'���������NL�蛞3)"�T�4��Ga��T>��$1ҧ�;(�UB�y�M`�\5��͎�T+��?��y���ѓ`y7��jN4�vp����fk6�{�?��?� �7���-�I���7�-�I��I@d"-w/�UG(�@��Dx.�^��)Iw���~��t��d�K�]���1��a5奭��Q!�~�sH���$Vi9��ϯ��
�S�A���K*^S]��s[��G]�{t�,���l&/��?N���mϡ!�m�����> 
!��T��6x�Kf��m����-;	g��&ޞ=���bd7��_��j���
�"<B�i��]bӷ��d���%��C(�!�|��i�`��_���B��ܤ�u�LV`܉�B�G��8f������(�g.?�q����Æ��1���h����ck�~s�ܐ�9�Y���<Kӝ��3I�:���:�l�R�W��N)zZ�LG���U�L�1�H�T&��#����~2�?��"���Lp�vb
��lW���e��s������t\Q�u���?�#밚# Soz�O���  �M��" ���c�UWr�Z�D7���K�8Eu��+-��1�иK�5�� q<����FZ��M�e����S�d���u�Is�a��L��pC�<*��|���6���7HU���T�ߵ��(�0U�#c�%��_꥾�gni� �,n��ݴ�+�������C�;ex5&ِ�+�h�yADM��G����kȿ4��SH^u/�)���*�Z,�&r��/�d`"�f��!�`&�$i��ˏ�Aǡ�Q&�M��˪2�6��Sc�*�+��}��+�V/������_TX�}	��?�!��}j3�<kU瘢��g#!���>��b�Ns�:�������::����q΀��L2~!���2 ��{��s:t��-����d�(��vA~��M��|h'Qޓ�)���@^
�GGQ����s٪ ����ض0�ԝ]4U��,~�'zEK�)r7��:ځT��1ǐ��� Pu�e' 	y�P��au�hVK��uk����:�xQ�V�5�e�:�S:���ܖU'E>U�0+��Tz���dL�Ł����6�Q�_��ui\>S�_k�~�ɛl!f�F*���92����0|c��@���k=`Q�2%�rkD�үB����0�3ቧБ;�4�Bjq��(�- zBj�ӏ���t$�9jwH�U
�2�9%��_	�t&���C�|�B_�[�4:��A=d��m�ǵ�9��lU�3ljSԿMzq��ǜ��G��cr?�m�tjj�`
KH�\�agJ�톈\Yv���n"�Q�rK��'�t�$�o����ۥ=9�Eq3W�A�&à����e�?���7�>o��׋�N���GgK��Ԯ1?���r=�0u��x�oy�/,�$u�G7�4r�粠f��cR��)��D�
����-37��G�I1���_WT�������Ls�u�u�.�0Gm׉��_x�7��K��\�ˋi�����)o��ɡ���Ǧ���N���(�=����bB!�ā�����vJ�� ���q��z��z� ��?(���9RQ�BtNj䑿�t>/������F#����*���4.e{��t�<r��g��
�0M�ĭ�I��ӯ��@�2+�/������3��G�K����C$8�	SH�)Y�]o@?�4Av��pO���Zt�.*A�D��C�3����$�m91��G��3�c�09{f����*sYʬށ�.�u�lw��5�_��&Q �'�<\��L> �=�\��<+��hH,�i�F:� ���5��-kO:F	ʫ�o��h��~�x�x��o���:/������c�ܙ	_����fq���Q�y�f�}fV#�P���f2�����C����h���x���\*�_�~?�5g����J�E���S��5k��_˹*��U�'�F�	$k?{PF2���C;꯴6�#A�V���H�S�$�R�FB��1+{<4Ź�R!�t�
�(�P)�˕��Ob����S�9@���s��l�i<2�i�0�'c/s#�����a+��&slK@�
Έ�lיI�0K�}�_!1�'@��`����	��9�i����/)/������!����G�$h�(���p�b�h�� ӈ	�(���;v�ӔB 'Vꅻ�	�����n��/Z;�ԉ����)D�]�	n��wqNE������O�l�2DC�QJ$�w�*�Y�PU4�5���}Mq���$N�u8��ݏ�x���������(X����yn��~�O�eП̜��!N�1�� �9U<~2n��Z���F"�E���WX��7���e�Ϯ]�e������������6���O�oqs ������]�K,�2�܄)�/Q&��}�q�Y���u�ᅧ��y���g\d�T�BgjY��)�V�;XWBΡ^�TIu DMcwX�<�ҼWo>�ό�� �Ī�[P�Qke<��B���挈8^��Ư_� ���t�s��>�<d��\�/Y���Gz�)�R�ک?E2�W��K̻��"f�\�����|Q	��׎��·�y�O��C�. �y]?+�Es���͵x�X�Jb�F���H�v�#`�8,l�2잞����3����&T��"y��n���Ya=6<���a��a�E�G)�z2c�������O�c����jZMT�sJ�/��g�_ƭ�f�
�#j������+��+2�K���G KhM�� f�v7�)�۫��������A0"B��Pl�(�p��$��s��a�$����Ŵ���;[UPl���5դ�\H���������̷c�w(�بp���~-�l��Г����9j�x��-��>)=������ܽ5��*��ٌ�B�F��8���/A������0��������T���苙��C�,�S��cPk�l� �6��C�ׅ���P$��NfT.M!/�a��^)�i舘�Ұ��X�ۅ��n~=p��E��P'�=��?;4�n%^�t{G�Y��X�@塬�=��9RMU�q� @#�`�P"�r�0(>S:g|d#����K���{��-�)�\Iw��W=�ZWX�	WrqV��C�r����@�ŷ���:�;��hP�ky�K}#��s��Jo���:,�s���'��"9 ���-���*���{� [�'�@m���1���Ú����LbEU�q�?�^Z-��v�t�4�k_g��j�.��F.Q���� _ܐ�P[���֬���ɫg�5���������=�p���Z���)���E�����uc�›J����Tw���9.�n�zr�;��%�T;�o\�X�%�"�~�fa7����f�f���0��yq1��|~������L�[+	v��Hf���P�K��|��OW� �N,8ꥈ��G�P�XmQ�D$w�)3��Y��x?v�7;&�e[�gÀEN���8��=@dT��B���,�)����|��Bʹ�#lB��Ӈ�����^qp	l/j�AI�����n$v�����3�|@�$�xw��I�&�79����e���r5��e�t�֘����p{yL{�]|zXWb�"�����νt@܃��("��Ŵ�ȴu���jep�����2:�(�5��C�]�LJ�h���G)��˄������55������ E}�x�qѐ��B�Z��USkYg_Ɩ�2���2Aa���͕��K�HAsan���Q�����	���*���A[�oe�HD�(p��4��A��i�6!��k
C3�ٳ�%��w�G0�����EWK�ż`�gB_�����˹����.\���s@�Ų��מ
���:���@#&d�#��������V�)��5ؙ�/ۚKa�qb��W�	�'��F�s�	�t�Ĵ0 �$ڌ-1����t�鳤�R�9��J��X��g��j�r�=����P�N�?A���zڌ���b�|��ZPL�~����w�������\�*�p��d�njOɒ�k8c,���.�>�[3�B#Q��J�
���ֲ�L��G��=�n뮌Y;P?c�:h��D
��?;�f鎇\�����}w��e������	V!6i�Q)cSu����U1^i��
Yk�&�p���y�
TU�����%>Յq"�y��kvi��ܬZ;�u�,zZjM�5��>)�NQ)���7�u��?+:�J�U�r��#�ǒa"�Z��J�%i���;*�� OGG{���ڨ6�Ϭ�(�Q�:��}a�
���5�J����Î[���/wVI�j�psf5ذu>��+�.Q�@���Ǟ���%�*��?��wc�/KQ��d�
���8��⦮��iC��Q����x�n�	�;M��!�6��-JX�"r�7N�����ܐ��@����{F�P�;}���B_u�2^���-�ȫ�Q2�޻��%�w����](W���2V�=�����j���<25+x�b
�� �����W*z��s�W{�H�`�&�F����B�Q�kT�Yzm�n�)蔨N"��8H�Ҝ���)f��6c;�)W���Ǐ����ꉣ��u��a֯�PM�&Te� p��EV<�rܔ��\Q	r�j��:,�!{���޴wo�\����D�
zCN�G �����#��.Ç�\`XI�)K�i'dr[JhHz}V��s�|� _�����EgW�-m!~�k���_�ӄ<w��<c��F	�\��M�H�������zQ�4�m�%��2};����  K��@�Ĥ����pt������QgYǏ_������c��q�A%���h�J�l��Q��	^�]��o�^�m;#o���l�F�X�cP��p�.�Q�G��$%��*g�'r��Z?&=��L����Ks�5#���8�^$Eىp����?��P�F6\2�ge�9���H]y�@���0N�M�hոh_,�j�_u�.W�5	����N�l���� �F���/�� "b=����Z,B��2 �iI5����A~���z�7wN�c����
d�C��]2a̯��}0�)�B()=>�7g�V�@�&�=nB�f�4��F{�Y�Pc$�)��~K��J�{�I�.�c�f�������|����Z"� �\���(~�&�S_'$]ܮ@�KU��,Coó�0R�.�@����Nɇ�����<nס5�Rƽ6�]���W%~3��`ZSHj"�j�.P��@~�o!����C�v�8�%?D���>L�Isx.Ei-�t�ev[�󅢣�����Id�\���|��ٳ┷��
8���=�������Yb�LxU�ո�ܑ/�|j6�f�E�6` �r�<�������in��w��P�۸c�u�7~�+�:iF�K��p`R�n4zl�5j4?�e��=�6��j"�3\���@�x���������������n$@ 1�3���u�>ӓ"��nh�)x׿Հ�F-��:���P>�k&Zb
4���g���	����'�c^sTAK�:rz�����(���<i�M/�dG�5Y��n�Ǐ�XTo����2ŵkς��J��!B2[,�3��>�&Zqv���iUa[����;~���B�������q���3%GD���ݲ+���ɮ�R���ok�7�-��Q-������x�%�s�G9`�';vL��H���S7B!j1�vs���9��sH��L+2c�R��]�R.k;��7���2�����(����=�r`� e�KtdP�A��y1��RM��/W!�͝�2�Y��>�V���퀨��#Z�%o^ɱ��t��йRK+pg׬w�	,�`����
��6j��y[�'NҶP�w}r�g�� �4cq�,T�PA��/逍�`h�&i�j�c���2����(��}Q͒�*�� W"R��;Ǎ�������P.�G>^FLb�x�@C��:�3��i�|�����K��;Ar��y!�t�S�{�"�1���(z&�,`��B
X7ɮX(�{+X�C+�r�Wz^	I��%�m��������b��]����7��mJu�1�.0-Y+�����G�I�ˊG��v�D��{���@3�X{��TF�1�$<���ʥ���NN�h��<ӟ&�
��>�f�;A�6<\"L>�Q�\����s�v45g�B��� ��tV��+L�20�\�ET��ФL囻 ������F�]�X3܍�X_�Q5�%D��Z&���07���\Q'��xl�����^���2j�\u�V�4h{#�X��1��g�b!Z��R�-��~m�4S�~!c��$�D���R�]0iB�a�k
@�k �îZ�����J�פ�.� y�C#F�W-K�o�@[�_�7f ����F�����f+0�4��������5?�xA���M+7>&{r�H���!.�8/�u偐���\T)��z�!&ޣ��)��MW�B),����n���b�yZ��u$�*�ʞ��r��v%�܍Q�ꋌ��m�'}K.�z�;LV�N�$��U�� �-�Q��u��;4��!)��o��kH�L�l��c���51J��@<��s������#3�L�[4�����Y�-�r~�M��*���^���	-�p:����\���nȼ�Kܲ�dv�Ϟ�<��W_�]̒�d[�//FaA?��|�Ƌ�ʒ`�_Ota�#�9j8�����{�\L�s�up���hE�I��������J��b�"i^�eu�9�:%D�5�_�#�8H���WR�/r�76S����#r$7��⾟��d��Aܧ��2	i-;<������i�5�����MK�G�g�yD�A� �b�,D�W��f^�V�6��]z�[T�AH�#C^��k=ڬ3%h]��+9�{C�秉�5�2ؐ}������c��ޒ�n.q�bw���m*%�ݱ�<U�;
�+��r��2�neo�U�9�����E��<��!,@��dS����@@p�Y��Q��R�C��������N�"����k�nn��Go{����:��Z�X���4"u�,�_��w��]" h 9اGٝ<��o�Q&�����!I�΄���d��^)[�m�0ˮ�±
v�����~����#U�ծ;]��lB��V��p�I��k�*󘞄s|�K�)D*�x���]�����`w�t�	�BQ�J�/@�rSW��Y�b`ɾҲ��r<�Y�F�	����u� ��fP����3��|�%) e��>������9���.�4��|q��2RʹR6�ٜJBK�Ůٶw�w��K��Qz�OR�����n�A��#Y�.7dUU/�*t�3k*b��d�a��V]ӎ�!��L�4��5<��g8��ɡH9����W��2�H�>��`�k��}ӊ?7�W�9���G����3��&�$�"�S�4cL�����(���������NM�K�zg���y�"��l{c��l�*�{�No�,/]!�!�X�߫ӟM���W�JOU������mi���z��!�~�A&��q;��pP��K͝u�;@uu��u*�{�|�Y���?��$����"$�㶏f��1��F$]$m��us���As]�Q�|�0�1������~\|���}=�:���ײ�O�>�<�{q=+�:�h�$|�}�VUS���z�T�����ͱ��7�`�S�"�$o�haXP��u���_(j�g���>xʷ���Я�S��9���Q{�4��Q�f��_)���I36�) �U嫑�D&�!ꞯ�<hsZ��	`-�z7@AhR��t��3]A�5�w~G)̉�;p�Y`�&�d<����F��I��̍-Äg&��g�����L���PN.��B_U���8KqK��֨�l�b(q�v�O�FS��䃽،�������
X�޳s,��BŔ�����?&��_�O���s�ݱ��+f�������N{8�{�p�b�F�A��1AhF�N-tg�V�%B_b�#���M>�&�`�Rx (���AQb9��i�h6���n����b�P��x����<?4�k	���X#MHO89��;�W��'L�CDE�n���W�l��3f�^5�EUw���;K��>j��2�jA�.�)��	�y���&��:��ƪ���8K%4ᅔr����Tsr�m�"��f���ry����t@d�%��/r8�jd�QB�Q�x�_}T���/f�\nb��Ic��H���.�s*N\qf�̻���z���MtZ��m� BH.�
Ja�\�B�SZO;������?����`:���f�n�%��yŗ^�M��P��5:[y
���M�A���nd�Jo�=a��%;��������9��]�z���B�;_��ׯ*�ywJ��),1�i�9v4���i����y�
�`�\���y�,ϐ_)>��Z���郊=M�^~8�x��)�ڴ��C�2��уu93d��[O�9H�bTh����/�$]~�H*v�Q-�k��,Z?��� R>�ix��(8n��j>*��p���F�d�~=����<�w+��@�wIT'�|/��j9Σp;k��U�U��+3�M��'��m<��1U@~��2��2�?��.fd(��� z5���t��qy{}�������[�#{UiHY����uҒ(ʑnGP��P,�F��1�I����(4��J�e[��X��q�;)����0P����=�-�[��d�B܍��:�p�T3p�P�ΨE�7U���B��Mg��/�-!y�6�.+	K��n��=ևzX$随���	���("z�֋/�Y��Ua\�X��.Ԗ�ʰH��g��C�zt��ZMs��V�9�a��=�2�Z|x���/8߈t�qQ`Z��ǨmFd5�`��3V�j:�$�`��iV{vNP����"Z(��`ԇ���ޤigs���qɯ�޶T	�B�ME@�J�;���lM�?�×��m�Z�u�ߤ��	p���j��.8QI��AQ��_I��ر�{��Q�Ԍ�gwE�
.$�^�����z�+���4�'�7���ϐ��P]��2�9�ῦi|=�F�с�P�,.�	���^T���҃��n�@M.i�$�j�v��2B�✠�(l���F��K��B�8V/N���a��*v�h)r��k��	/v�'�|��!?s��E�̙�9�u?��q�jD�l�@��˲63y|��ܣe��t-sS�*J�c�J4���+|�5��v��
��o�0=8c��������߯���q<��>R&��gT�'B�sP0M��"�2~2��$��3�%��G&	M3W�����z���=Q{�-O�l�C�Ӣs�:#�lsj?kYx-k,9�"u`���m��!��P�w�c��:��R��k%�W��Ö��\�������ۆ�h�y*u2�0�o%�/ᘹ��z�)�N�v<;VV�\� ��Ǆ��G3��Ã�Z�ڨ׼|��W�E5���^���o2!�Z���L�58��v���*�ꨆ�k���}l_�"����^��.��_�%PMA��t[�oJ.������R~��]tC�M"Qv%�j�/��S�7�J��X�7�V�M��$ � �s�v�DY& O�)I����v~�X�13ڭ�����f�Ŏā�XZ�Z�bV��ށ�'�p:�čx��n���H�S#������.;_[ೣ�
��������	�\��L�0F쥻���p��@��J!��@*lQ��K=�Ŝ	w�ϋt�b��Q[
��y�'w��:�����!^qp�jN�Ea&g�4��ضÁ@O=��"�
��)�Chd��A�,r�٧F:��-71fw�1<����;��BY�@T�����c̎���/M)�~�����DC�bUZ�Tv��%��p'��a��1�U#�XL�������:���0|��D�5(z D���bp�����W��0����Pep3d#_V����>j�dk��3[�j��a�|��{����6���Y.aNw �NO�!���:zxhp��?xO�6��ç��`�i8l�պ�[<W���^�=��͍5�8�K�eSL��^�&#�y��P��ʽп�̣D��t\3Aj9��	�YJ�Io,��'-`Q�],��Yl.OTݕ��� ����C��LOSR$��^20/���|X�ۮ�ds
��#�¥���������ꒈ��l�<{���-q|Wz<`����G��RT�}���bo	�V�l/ ��4�e""�N?�j;�U"Q�����^���5kv�oK���o��@>�>�De����,�T�������l4T g����4� 2��n{uQn�y ��_1�`���*��፧�Yr��M�,�v�W2|�Q�z����x�8�~�?o�O��A,�ȫqQn���5਌���q���v�j�:G���/��q��,̘�*Ĩq�����9���O��b����/�]���J��CeyYA��ݼh�� Aq�	�U�*�#�\�Q�y��u�{wr��gH���S�vu�q�[��R��*�\���:u-�OG�'"���?�3�*>���Q,0t��R���0r�_�A�����!u�xl�Bā��S����Ϯq�aKe���h�����vnX�"=�4�m���	Ej6D��T#�j7�;����7�+�$�X��Jb���b������p�4�_�[X'�ߠ��{�^�S�vP:;�U^<�T+x;�?t�OK�4m@���'���7����޳k�n��:�\p3�O�'��R�fݓ/`W�+}�6����܊R��(�k�]�� 3R�>�؇�|��"l�R�)I�Hjj�b��i��ȗ�Ў0�%"ͮc;���JEcC
����*�"����M�o;�eZ����1+��dG6�F���b��cR�~��ҷ�k�(��	��2oە���,8떞Ik�f���-T��VϤ��z��N~[K�̬�{r�>U3�Ǌ��Mtޖ=Ӎ�8�!�>��!�BN�� �chf����e㓩�IYU�1��#J���Xb�`tS\Bd3>u!Eh�R��J	K��MR#:�i���0��ǐ,[�ۓ��^�fםЇ���� �Qݛ@��	���-T��|���X�,��q����R��)��@��P#KBW��⬂o���U�۸��L�T���僽�?��V�he�/�H�s'�f4�:<�{���>�� ���K�R����T��{6��l���mPTX3�`��|��`�%�T��dNv�I��o,e�e�r�!��< 3�x�p��Z(l���������Ih�qFh���«�+���ͯ)�nXߎ:^Dv
U{n>O/�%�Mx�� G�:�_`V/#��cC%��-�s6VU�,��U��x�����
.�e��Q�c���C���;��R�����Dۓ��#��i?��&LrCtG*ic���R	pQ�\P �
�\J��*�A@.��̷6�����p4*1�j�ȉ��h�����!���/e�//nUX}�<�ӟ�-\8"$���$n�xs�b�7���5HhM��b6���+i�_k�S;�J-dw��{p��p/�G�.z�J������[ˇ�J��2�`+��
��`!�Nխ��De��˅Ӎlc��C-g�i��?5�M��!�)�vDJ�����ۭ@��~�>�L������H(f*㯗��ѪF
[��F}�dԑ ���s%��V����EUG��-���[�E��9s�`����u��i�$M���PSQ.WA#<���Ɲ�2n�����!����d#��{�!J�h�^NC��S~��B,���s���M���Ǫ��
�"�2�1���O5<4���_7�����g�mo���;v$���U�FFK �uهdC��J�_9�Z��	��e�e��U����Ua����cH��0���~�{V�o�5^��ߓ7`�@�K�-Ui��>��:������H��|���9PD8'2�����[R����O�۵���H���#�W�Yl3�F�N���9N_rrk��/�U�s�ZW{�#tCs�.Q��FL�`+<To� �y���Pyrzj@#$��vPB���c��ɝ�bQ�^F&���9.׼�U�����P��
��d���W�߄����k�y��U�]@������pM�́d���5�>^��U�n�����H�&�UB�f/%�E�I����K�fVE�u�i�5��@-�V�0����.���1ˈbc�%�"K8�r���� �oj�[J�＿ׄ����1|��413b���,�a:�^#��~,�h������#�cԊ�鐿R�p��޹��!��N&��x��Ȍ���n���"�� *u/�/$�ߜكE�Wu��Q�u�Ʌ���zey��L�
_�r�[�o(ѩ�SSL�Z/y/冉g�f�4j�tIի��Z�o�\hVT@�]	m��Cw8�{\�]���*�N@U�J�܈���'U.�L�V�H������dǣcF��~~��Y�נ��Py!.�F9�V3���Iu�L�e)L�V%�=�x*v؈�|�i���x��_�̇\X*��Z��"�ؑ_��ν��ϰF?�+�	x`��~��&��u�b�̯^@��y�����e���N�2�YO�({���W~b	����~��u�����!�",�8K�1W��ٓN�25�_�]Bf/�-�y�f�=�EX����혭��n"'��5�(�8�As"�,�e�Ү(��JoƂ�m5���CK5�;V�_�+��K�Ac#��)#��~�n#������]�7l�D�	��E�[(��"2��s�T>GK�4o������L�(�����g��?���)��mLҿ_�QVX|�_fZ4�~���`<��r?_u��2k�c�;��mf��	>q���6��b+_C�{Y���럺�u���`ՒdF����ƒ8LL�Oc�+�Gէ�fH�k/��7	1�h�qB��U�z$���9�Ht����CF	�"ˠ��	��]��Qp�������o!��N��G�����	�%��Sx/�D,�<�W���� o}�Z�S0dd�f����q����Ǆ����*��̾���n����d76Խ��������r��%l�RR[��8r�u��F	☊6�p��F�e����}� [z��q9�f�3�޾�ފ�{�S�Y7�lz�U~�6��]�uZ-��ǧ���!��M}�+���(Ρ���<x�˺E��;�ﯜ�j��Q��l���C�ҙ.¦������l~�SF{�N���f�a.��S����6j;�8G~C��QA�_a����Τ������5m`�$_���clL�E�iX��&f<ڦ<Cd�!>(�,M2���ȝ�"�[�?��i�����9	[֫��P&�cL䮠�<���~*�x�%vr[����0�� �ߗ����@|x���9�<eo�ǖ�����zi^�JQ�T���K;�����V�ѫ���ѵ?1����eC�u_�t�N�ܻY �2�Y�;36?�R<�<3�,}�6\$�Jj�V����MJ�!eo��Fqr���2�pc �R�K���|�ȹ�I�p>��g���f�@�$��Nِ�8ì&A;t���l����