��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�KW�UHս����fP��nIw@��Fn�~�}��w�{���ڽR������_^�p��1��q�ڪ,�S鄄(I��jx}I�����y�"˜idW\��9� ����l/8�g�UB�Ə�7��s���#���&��4�Ũ�/�85FLHE�t�)"!�}�F����L�AfY��I��I�I�(�I"u����~�t����_�ʶ`�R漖��-twz�S0����R�	ōU�ّ@߃g��Ϊ���|4±��P�Ak�gvQÅP1��p����4����=�_��j�l8�5�\��6xc�����z"�����|���!톼[����g>o���;��W�yM���M-.�E��4��r��ve<j9x�hL_�
��Y��O��R1R�����~���׀���u�ަ��b�,$���}�C6� ����S�w&�A��h�3��,9����KYo�[�b�E��$�`��t*��>6�� �ć~�����k��Pe�����	�M�K�����~�*�ʆ-P�ss�;��>8�[O��Ǣ���Z���+��-DY�����r�;XdR�$�dQ����UI2U�}>@7S�6��Ăm�Oև�,���3B'����1o
�[~��MG��+8�K�]�ߔ>j1+�O��->I�k�y�u$�+S,,�M�kq�j������W#T�'�I͏��A����<�����t� �K#?�zz�{���@���1pJ��}���jdza�
���R	�]*n_�JT3��z@r��W��le�z�e^��V,�v=��$�-���zɧj�0C`z��[[b!{�E�$�:���<�����IB+*������ŭf�<Iݾ����������$dE�M�wO�}ĿXťq隬�z�0l�e��n�����B.�&�j�[0E�	IT8�����n%�ˎ�	-�O�"��ގԚ��z� şy��m+���P��n}���C�\KM�DoK�W��'~F)85m-.�_83]e�eA�'��Q��i�vL�Ƈ;���P�#�3簿+�I2���!���p�u�N��$p;�.�f�5QB5XMs�(�K.�ن�%��f]�ia�f�M���d>]a�q ���l���\��������l��Ƿ��p�b|}����1sxJ˞���$��������p�i}��� |���^H�p/]@c��T�W�0���:5I89�jū���� <^���g���qB��w�qE���6ױ~��T$�~=��K��̓��KF)�XIg�x
���f�p�r�;B��(�;�Ę�$m ��_�&<0�G�ݦ#�X?�W��L�t��{���lJ��+I0�
�m(�e�v耪]���;�\���1�˄��WF3��+8�u����U�=�[/�o]��$d�x�T���4c�Q�,0���u������l���ɫU���'J����;��: �ۇ�O�����I�#_�T�|+˳�L�n}���eX����>�5n�O��)��'�^�
�������4d�.�(��"보��#f&�X�2�ȗ+�Y0���)�Z��ق?̅�h�Ӊ�|�(���A��,�N�2I��lմo
���o�f�dC�Z��/m��!���?5���'��0"�ʄ����󱦎1���Zʶ�J�#�=�3��J�4�Q��>��n���J�X��1�˕��i$�9k];�7�[��C�WE�nbD+MX�����^���t�9>y��g�� ˯��">�f�
ֽ�b->��K@��Y�U�����3-�=I�*���:�V�O;tJ��.�i;Z�%HrlnXf�!���,�%OA#z#�d4O�"G������,�g+�Z`�#��"��:�a+R�=�>�jc����CmP��#1�y��g�x�ς�o�w�I��C4J�u� ܏&�!h���m���g>�,��1�`�!pK���7!��{�o�E��g,٫,�g�ݏ�b*v�\9x�ݽ>��W��U%��v���^�ֺdd���X����١Q�Rǁƃ=��ߋ����6
��A�WaPU-����О��{ _Y>�5�p�����ua�2Vr:���������j�Y=&Τ$���9-p�j}}�j�ޣ�����OK����� b�co� ����5%1b��[�����
JߛW%b�Fqݢ>�O���O�:Նd���F����5>�@!��x
-)��������V��	8��;��v����ݩ?�Nk����6,�:h���˘J��Oelq��ϣ����jY;ܢE�t_oz�zzv	�tF���jl%��=��I�N����Eih#���@g�M����|$��'6�o��.J'#MD����!3�����9��(gZ6�]uy}�~����w}hs|6C��'i9'�F�is*;�ʄ��#h	?�~��\��$�H���A�".IL =�oD��;e��[Gw2pk9�������ݞel���;�Ҿ�}$k_��'��x��Bh&��O�#0�pנ����}�Sa;t )���}�����}��i�a�X�JE���,�-��&�����1�2��r�$b���E���V�N���=p��S��9E�&�X�Gs%>�"<��=>�郄i^�[��)w5�J�K�%�p��w���qn�\�\�A�.��2܃����_7��od�?'>���K5W��N/ec���c+\�)O�S
T��y�H10���G�g�L��B�|�._s�e.�]= Kq+mh��?d�qe�BCU��%��؀�vC*u=٬���"�)�g�����l�ףY��H�����&M�xh�9�/�E`���}�:��9�=���ؠ� �!-U%wJz
�t�� �
�����i��ad�OFH2��4EBl�$t���C@8Z�K� -��&�I�N�-L�S�-�S�H���\$H��IQ���`�"@��R�Ŝ{8��ԠⲚ���g���帽=���)|�*Ɓ�6��r�T��\㈆��DĄ���1�ꇑݿzT���T~�t�)��{UrN��Z�#�;iD���������B���I�6$�ș�K��mK�/��f\����S8r�:�̌��?A�D�"�͈�R���x~|�����WV�@2�@��S�K��#;�օ�ai��0˨���	%f�s$�ܮ�$@w��z�}Ew�d����c�	��>սB�R�I�KY:U��0!7�%P=�n��x����eH���GR�L�� �gU/,��.)��h#T��G;h�r[�y�6�6:�dc�j���&������)W�WXn�rC�2�Ȅ�׈Iά���!r /1��;�|)M���+(�6��9�0����R}��<��/$�� o���X�uon����x0Bb#���R�F�j���l&r�z2?�Y�?�KK�Z��v�2(NѼ�Nf@8�p$�رQ�����u������-��ߥ�"��a)Ğ���\���2��#y��!D��L���E'�0���*]����W��ѻ�'����.�99��?�r���Wx��=���|�{+�W�<JN�ȸ�������1�_���43f��@���������_�$g�#f'�)���,u����2����/� ٹ���\�OQ��+Yi������Z���2W�����3����'����Ogu��t~�[��������66���Pv=kQ!�	��Xb*�;�H���^	􈨓SB�4�K3�6��I����I9�k3���Q�/��+�������7${&�e����Up��	�����@�P-;�G���U
���ZPR~ք�����fE��J����N�]�q]7C(hUw��;D�]���?!�W�"诘�u>Q0�L�Hy��D}p͠ �����Zv��ʉ�ֺۭG�n��4�~�] (B*����d�F�6A� q�D@��#eOđ4n �1�!���9@��d	��K����*���9>� L�U��`��́�]%|�L �Q"Ptn)�OaSl�J���^:��赤�����l�H���++17<�]dJ��F��0�7���7�:�3����v���O���;k;�?Y�0'��3^x�+|AT����c��M7pr�	��ح�F��t�~��8kqPFaW왦�J-������,���UT{�Ic.D���V�RyE�|R ��=2oe�/���J���~N3+��&*d�,�ư�I�J�|�(�(��2��k� �W���u�K��g��4�4�­�g>$��C������{���7�bg�9s�Xg�qR�	$9��3Χ�K�a��g��������ߝ[Z�|Lj�0U����U�-�2��~p���X��o���<�:ʰq����',n��o��U/����gim5�b�|s���Y)��>2k�^������H�C��`Dbh�k{�������Z�Vh�7LΝ��j`)�i4|>�ܽ��>�����i{	Q|i*=�-����&�8U!�<��C��D9��;?�����:&��U���<�	)�G1���|U�\��I����Ŧ'!�����i�UT)lZ|z�b�e�0j(�_�..�H]�@���r`�Y���Pk����å�di z��^s��q�T���3��Z�Ϣ��%������w���uV���A��G�����-��.���^
�C�6�Է$$�C���@�0ߛR�Y��]c���j+�ğ�F|6$q��2t�p�j��D>�(;�	E�ks�� j�h��;^t{9��^��,;H�t�)g�t�^�y��_ �C���i��N!(1�xl��_/`�	#A� x����8a]X��c�y߮:Y���	&S=�10})Q>}�b�I���,B��P�P�lPD�6)��}�g�R�Ӎy����$��Z6Vy�rH���H�{�����#�Zg�W��b���b;���įƺs���3�Rn/i��Y�k�� ���#\c�-�2y���G�q��K�	s�O8�IG�q��YfS�9'��hF�9�Ts�A��	8��g�ö``(oҽ�� 5�;������3B�~dB/��+HQ�℩�����
�HTE���*6�q{�C*�%i�!��;�X�{+���J_�6�R�ϖ�ǈdT��=�ٸ*#^қhx��3�м�F��g�f�2?�p
���N���w]��l��,b�e_��.T�����ǢP��h�O����0h�k���A�����>;O���N��e5&HU�O��s�4��ĥm���7(D>Pg]�Z^�ח�ΡK�:��3�):�jW�N��]�E�^��<_�L�_1ľd�N�����-q��O�|]�q' \
��"�p��+rH���{��Uw�YKJ���x[��6SP�x�^�uY���@s��ā�vA�v8�-?A:�1�����fF��Үue�@Q��F����9��۟������Kj<��,�x�[���Mh�y0�*5�:' 1�`�t���Q��jb��6O�Μ���{j�����O�e
 ����W�,�<�%̫T�gP�+Y;oe�(�t�t������/wV�3G�*�g�
�^9�^F%���E�/1���j9� ���d��ebz�Μq�e�>Lk��E��q��6�t0���}~>c!߿�G\�}2裠�Eޫ��׽��/S:/���2S���j�'�p|��B���8�4<�$����ٳ]�[7��Uj߬h�M����S��q��|�2��]���=x���C�"T��ѩ����}�(��C�V	���$��~��X|���z�=<7�<S��:�]��~��F�}U�jq�2�h�o^|����J��6�K���NG0uL�,Xc��LY�O��.]T����JVx5��BE���r�@�P4��Z��y����qb�������������e���ww��q,d|�_v�e��'sJS:�n-���C�v��Nw���xs�ī�%;L}��[��
���%L�L+����������Z�i�{@��<=����\�t���x/� )ȣ�:Y�(�n~9;��%�q�fʲ�!��L�������C��$|�z	�����$����b�W씥��fh���}���򴻂���F�&�6x�[���P<L<�P��+C��2�1���.2�JF���[����F��+2��:�k�O�t�Z02��k�*�����Ja�䕖�~ 8ƭ&wq�yY��\$E�� �b�'�q�̝yܲH�n�o�GxQ�u8o���B � �[��ۋ��r�=�]���X�����u���B���b���]ԕ2���j�?h�`�����X�Nb�m��c�OTs��M�͹�����-<�'`�"c������6k�̨A6"����E��ϳ�rS^+���� v���,ȥ2�"���G��m�O�o���A�2���d	����i��):֯�n�s�B�1����s��S?��!�
Ir.*aA-��DV�؅����<�C���	��Ch�ҕJ���<�KT|%��h/a�ؗ���K���V?�+ajQ?�ɷ���4�s_�'6�G�����1���W��v2��J̗K��5u���o	#@x�F�.ПN�Q��ߘ�r>e�,t�0�
��\:G���nnF-��� 6����eC�skƼ
(�&�[�̴p��$;u�u&��5�6��N��q<g?�Μ!(ƀ	C�pEe�����#�pm�~%d'�lE%�)�#T�-���}~�sЛ�y�Қ��>�
��Ggf�[��B� �;k�ϮR�ʑ;3�m�Uq~]6H.|�Y��*G�֣�L����8k|��DX��>	 ڍ&����h�~�о�`홨G�@��3��:#�/��4Tx)��W��T3xݳ4!�,յ�A��*��y_���:	�wmt��j�q��_�}���C�	B�T Vl!�fX���=$3�F�\[0�sS㜛�!�1�>�	vQ����}>Y�D�ӏZ��݃�!#��M���liP!��Igkd�/.��tم�p����)x���F�wT��"�VvWfX:�)Fn����+#�=��<��"U"Y*˳d4_^m#Pި�1d��9�pP$�/hï1�~�@��{iq����;�ܞ�󘶺'E�i9���̆�,5�T݀��#���'�_��\[�����i�����8���x��:U�FMa��Q�P޴��n�m?�ж�$Ж�]�p�b0���~5bk���FQl/]��)�z�.5��w,�Ǵ0�UӼ���Z�=�Xf�J�
lc|C��nA�^�lYkM34���Hla-�,`���UO�I���G�����Ǚچ��*���.2���.����W����~jq<��2 |�(��Q�����be�^���`Y$[X/����`�.���������A=BJLjjaXQ\�@�\�����w��n�U
qw�ħ{j1�k��^J^k؄�t
^��"��_m��$��7��K��%�b���=���71�S�T\\�IR!�.$A
������d�a��X,">��}I:UHp�_G/v �1�Y�^n2��G�������&�_���(��Dp�y'<�t3�lh�}-�@�G��zAA�m��Љ��kdx��� P̊���C���|���o��� �wrp9���s��\% ���=B=~)_�M�s�Q�1�0�=0���/ip��ǂ���
��3L��{��"�L�{`M�a��V졓7�f9����`�E��g��d�	
gt��|��˭kA�*U�#��S�=�3h�+b�C{0+��?�=�M��rg���7��=y�L��b`���Dn��Qs�#����k�)�#�+�ͥ�Ul4��ķɏ��)��hܽo�^��X���l�Vw��X3���&)f��D_sU�:��S�k�Q�$���@FwӠNzIf�\;� ���x'��"7�΢czٺ���������������ْ+,�:y�f��:��	*q>Av�z]�c�������ͯ)gll0���s�9�.�H�����w��_������Ȇ4��lo[u/�B]�h��G����0��9D�������E�X�v�w�������:�buo�����Ke]�v�)�\.�o�;��\Q.���W}����X��:販/ƞj.��`ĵ�#�q8�j�v)C>�~qM ?%�F��2V�3���w��g�C!}�c��o��QT[�����˜1�u�T���I+	b�A�]�a����fh���
V�<�k!e�	0bw ��6����6b5�MZ,��_\�M��T������_l�S)���nk�04 gl��>��s{8��˪Y���ܐ�(Q�x�������$>�x��{�>J��'���n]��NzZn�[�ʫTƀ)�T[�n��am�@����G�Ȭ���x���
��0d/������r抶�i�@'E)܊��������2�e�ߨ�I�������#�|���,4-�	΁�����	}�l�)�X��,��0��e���'����Qb��<<��<�I�( *�n���pW���4(gQ7�1d�b��R>yx�h%�9��YM��R���]H ����p�'��b�h'ג]���`Z�^(bC�h0��%�����ү��*	7:X�m�BǴ��Ivͨ5e�W���𚶉��#�=�ϝS���vx�¬���e�~<��2�K��#�E�E/yI]�U@�)Wpnc�e	����l���}�m#��k-�TG�rm��=�q��:� n�ݳ��ːH��F4�<��gͬ5A�7�:W�i-����0F���F�����O��=S�V�^�o��971̽ޜ`o%���'�9�u���@u�W�S�^�T�/�� ݝ��#�+�����J����H��K����+�fU����1�����iPs՚ }\�٬������*QZY(���(��h��-AlC�"��am]��`�h��I,w /C��Z�e�����~����ō� �gf-�0����C���	�`���Wz�t⸢���3�2?g"'�������P �9�ίZ�D:�n���}z�@ԯA�G�,�u4������¥�M�xk����c���J�?�G���?�I,���uoZ֜W�·��A�H�E��8)�$��S�/j��g��$!|�����o�2lNy���iDi����R8f~�x!.�[Xp�ֽ|4Ϫ�^�kr��y�I�d��iy��Ջ��U� 3�dMg+�����t��Fx��|��:\�T�,kh�����6�������DF��:��J
���+`��SJ��Z����O~��o#�-SK/��t>2�jƐJ�^w�?K�p8U�	-5�HH�'���U�]�+��<Ï:I'�Ħ��Y����Ō��@�4��<���G������[G�����!_�8�<q��_,����a��N5h���0���%�7'��B��t�B����u�K�$��Q��L���@=��`,���+!���3�������E:�.}̑���^�G�_���m �>��/�S�J�_���`D�i��~��w2 �a�q�vΫ��V�W*Cu���kn�W�V�0M�k&�UO��`�&U�9@赫��#T���u9���UzSq��	��!��$e`wG޲���Wٱ�p�Sn��^���X���L��O�^�/�	q&p}���%+���V���@��/jT_��~��H	x��T�����fE[�n���=e��Щ���([��	'�y����ŗj+h�᱉���.Ł̔��:w��D{�:�/���m�gl��J9���:�����F%)�l��=���ZY��C ��_���䤪ly�3k�hY!��ڛ8C�C�`g7�O)u'O�ړ��H^�Oo����ؚ�e\R���FE�q���d��P �����d��6&���,�N��Ӥ��O�l�z�sV�f��xo^�[�� ��K(yVr�H4$�[1 b��B'k��{�B�e��k�Q{��	�f�����y�YU�EG�*ݧ���Hq?m���	�ܢ9#uH��,�=�J`"M����l��>�+m~���櫃 E/0Ŕ_O=Sq�K%�ՃI��h��ڮ�J�Q��g�g�5�4�<t���['��<�V��+��<8^�~���H�)��=�YbYЖܐg����^��Lk����u�Ќ)�Ƚ%��Y�y�E���cI$s�hf��.[���,R�0O���)iE��JT��)�!�YE�o؈�x}�Z[�Z���U���i�F\2�Zm�?6�Њ�úKt�1�Ԑ�������5P��s~ ۗ %��g�a�<���4�������{i���LX�����xR��۴XQr�3�
k���[�ف�V��3�.q���f�C�8hV���d* 3ݎjN�w�bc||�k.X�L ��f~�E+hЄk4Ӌ"���x����u^�b�w�rFW7k����ф6��
�@�s�\�iw����ϘĶ��o�[I>�sN���eC핇�e�x� ?�V�k Z�8ĢD��[��K�:ڸ�/��;�س����>�����`��o�m�L�������h��O�n
М1毶`&�:Su��?8�+�K5��}'`Ә�.�{<��z�P~���,ɚ�������_L�M(�cͲ���́��(����.P`����?݁u�qW�G��L��2�U@����T��9q�i��7ÊԽ�Kb���ӫ��(վ2ǈ�ʎh"��M�6	d��}�Ts���JJۧ� DBB��`�`^���v�.��^F�&�X��V�FG�r��:�f�����#�#��*\m���D ������ߗ�s�x��Ѿ�v�x{:l�p��Fi�˫1�d���OS.��)flP�f� �Ly������J�Xx<�&=h���I�R2Z��E��]{�c��f�.�U`YI��0ub�ǲ�笣y�$���EH�d|��R�UyiQ�;eҰ�H��zb����# f	G��_~<�]_�m��/�1���t#9��x᷊e�0�{0����1͙����|a28I{����5,�8#4Q<@$ �ћ}L"|�U'}�O����V$�4��d��/��f|���J�8?2sA%O��|���EK���q�٭��Ї(?P��nk�`{�T)^R��N ��.8@.�Q�����ɐ�g�:�r����=S��<)��L��dS�b1ʱ�0�4�-�V����IS�G^�x�Z��|�|n�t�-�X��B9)|t��D������L�kc0��m���y�z l�/=]	(*G�󍬘x$_�:��ܙ o?!�|>�~�;g�0���������<���_ $������>"����=c����u�>��^D^�V49�*�	�%�rݝ�e*QB����,�*Y��&�3���U���'W4i�w�p���y `n'(�R�l������#��*��@���Fx$��Vw7&�������ԙ(�ߤm!����6�T�N;oRz��9B,���w�g��� �"��jfK����*���r>f&�ђ��8P;���l�o�F�Ul�9�cG.U����1�7��շ{�^���:k*�������j�|h�V��dZ�ωWG�O�l�U^r�@)��i��ش,�f
��i����3E�)xJ~������-���`�֨�yǌR<�����Λ�[��{�wD�?g��22Q���o���UD}�� !}W�*�۶�!i�/���zݍ�����LMun. '2a<ц�0їM����Z��03��N�W������7�+��oZ��U��:��%a�Ñ���� �[7��{�i4d��;G�S߹���ta
�ߌ���%u,f�ߊ�?؎ E�%DSE"�[:�/}_�aY�D����2O��Ӭ�]z����t��^)���7C���X�a��c��ͪnG&��jk.��̋�,�,�Q�yӰ��1n���Ww�PJe�Y]k�I�9k*H` _�U��r��%~����Ɩ��đ8��aB�AJ�%\�sZ�X]I2ycD��6~����8��"���l�c3�#*]���<ށ�]�'A-�%����-��T&�-����q	"Z�#�����~�c�0G�NSBc��3��8ҾχM��������|k����ŭr����M��v�����{��[nETX#����(|7����=IQ.�%�)������>��P@d;52Y�DjU�"V�к��� �U�J^;!����u���6��ED�`ez�!¾���Our���s��+GAbrVS�o{�R���B�U[�ݺ��^�	i"�z�n}>�g�;�ڃQb΀7K_�9�z�_)�P�Dk+�H��׵A	��k��.��e��AfNu�4�����̣��^�r�ݼ�0
��嵦彑�J:9O&�A�QI�x�b�:�{2�.�=����0����Q��Θ���/�{ED�^�G�;(6F�Abﮔ�N��1I~�vW>�MU���ZE�x|."GT�G�U5��mR�|� l�|��T����,2ھR�Z� |Q����!����{&x�<������d�0�UR?i��P)�Go"(� C/Ԩ�
�Qc��zS���#Au:�wl��5g	��z�Tl�*�6�V�if(u���iŖO���pZ�o�b�HaA;3e��(���b�:�
Q�ڦ��3ƣ��Ѧs�qӹ=�P�˔��`���&(Ζs^!�R���uQL��z�!��{=�1/�9:�"S���ܙ��j�S�G/�]�w ��I+=PR����;��J�ґ��$$�ɺ+f��D&i	|�
��uz�j���h8�`�)��}�ɇ�ɕ���O
W�
i_-��58${UW����QC���(y�I�ؘ)˻�XS&[��g�O53p�,g��2�l|����s��AJ����]�h!�ޓ�� �ѡ�>�h��� N���֝�m��Qq�ן�XA)A���ӟ؜]Y�X��K߿2C+Dό��kb�.�e��b��#5�
I�?���3������MM��3����Ɩ�l�ֳ����L��rc��Ba�ž�ɹ�/�@�WG�T�g��� � �2	�HA��2��"~���9���Ϝ�^�՘V�t�!������-8��!V	@D��3.�s�h����̯�i�$�J�6KmW8�q�)��d\9��m�CѾ��w�����ä'W�}�TZ�?O���ޔ�­[ި�A�%|�pl�J�0���9�-`iAM8��&(%H`m��iuV/�ݖ,�P	�b�v�go#��|N��k�~̱KcW�Ɏ=�'��v0�����昞�G
�#�\���w�Y��B�
��ܒ��.0���}��ޡg�|]�#�z��'�UBeL�NP���~Q'���"IJjq?V����]4�Hqg�v��r�'�S�^Gf�0��=�}�ތr�}���]�H�q3�/|�
�Q� �&�>�s�'�*��9�A�Pݙ�b�u��[>��f������!��v	�}p�4W�z�=��F�W�:��;�z���(�0�5��vm6ڴu�����o�pjct)̐Ke��5�w�/��,(����F p.%��`?ч�a�J�6����Aq���ad��)_�8�X.C��w���ĶZ�8`9�M\lſiI�Ʊ:��ӡ��$ȊQ����/Q���nNԥD*M���s�/���W�i�й7I�;GB1�h��ƌ��.(�0��\�WpӳR�}��u>�fң���펲�x�q���J"	;�H�
v{_���~S�j�eG��O����gǌ;3%��A�#�����m�8�{؋Y�~+Tǰ��(�^*�Ӧ!�XT��Oا�A?��d���G�o�9�bPeb'[s���F�)����m�_^!�k\#�:���+:��f�A~�3�\{љ'���*��j�d�~;t�y)@M�
�N�W찝9�rY�P4$�uh"���<�o�Qx��J�VغvE#��&���_�μQ�����J�a�3�GC�*&���k��oh��{�g:S�b*ru6�m��W���N3-�޴ϠN�爍-�lY�-�]�L!/cW�T(�ȳ��V�����67��*��b�GR��Р�e�"(�9҅�2.���n̹l1G��b�&7������1�����$s�}��p�=��U�?�>[��^�)ӭT��%^R�iJ�4:&�2)����cQ�[���;Ө�1�����=MRF��ז�y��ݚ�Ҩ�&���󰝗p���dO�;	�;�7�@`/��<��)��Oخc�$\I���K-ʊK�YyMk���N%��z���)���Hɘ���+]\��G�:)e��Ҵ��g�BI�dx�7�Y(�@��n�]ջ¥��M�|�5(���>-F�a��0}�Қ�7�[��7et�U�u�{�)M0�[K���
u�>qH�W^�9lTwb@r�Zb7P�DJPXz�X1p?2�Y������mt�m�W��/I��]m����F�F��\U+���M�z����>+�~Lҧأ�;�豪�z���&�N�B���v��BC��knq�|UM�C���8nM��Y��O$WQ���;��YN�A��1�1ǦF��ӧTL��M�Ű�,��L�c!�Ӑ� �F
�&1��DeΠp�9N�c����p���0v�<�OU�H�a��j�����r�򑞞|�157e{�էC5��~���>�� �i�"��.��X�{�ݞ8�#��+O8m��e�1���a8p�i1i�pQ�U��1��,EY���5\���&7}�0جbT[�(HY�&�!7���{M�v��5�f�va�lK��s�ˆ:�9JS��i�y��@)��g��+�w�Y�~�=�*���~)@�z�/z�OOV(�C'�L��:� ��}��ݢm(e�dN%��S�����O߅�t��x'pU�؜��nm�5%39E�d��?-�RsHM+A���-`�� T�S����e�}p�wA�_F�p4�Y�oY=�!r�q/SVSQ,���C�|��c�\��^i#�-n�� �
��7��&1�H�<Gw���p�-�^ƚG%��A��/ؽ��7�B�sD,C�1�"뽘)��}� ���~��}�}�����o�DtK���#GL�	g������U�~�J/��kU�9�X;O��<�o��>o�rZC_�3d�E �@�������|�H�k��)�����X�-<qC7��^��3�L9�g-c�8�YKW*o��]{�SyP~b���/���yG���IΡΪbV�-�IOB�شx�i�S��-�p?B8�3��U�
�d<<�9�}����l�+�<����@r�ä8�_���J�����Β��'���|c�U��A��kKap"�m:�!9x]ƭT���2��)�i!H~�YuS�}�'K����N�%l�� �8)��;��A1�v��eX`��]����6�޵ٜ����@*�؟��E�%�-`���j��
����]��b��S�o�_���&IĐm���T�����ҝ9��'�b�H�>�*[:iU��o2��eC����&|������f�ڴ���?�t�;U6�C�B|C�:8�1E���I��@�ə�s�:�-��k
� ��� &��}��>Pz�N\�]v�P�I��*��Wnٞ��X�Q�,[5e�a���LJ9:F���D*4u�b^�b.ׁ)*���c�83�3��]��#`���MY�TCG��!��c��,�AV^�b�Qj ��BxI
���}��ܧ'�0i�>�9ӧ��fM	��S��\���beN�6L:�һ|!]�hX������hY�4a��qΞa�	��s���լbMKF�
W� &�4��|������s7ǔB�5	�����g���R\Q&/Q3
Sd>�+O�����9>���=4-��.�p�������l�jV�:Q�<��c+D��m����Z�y֬)�a�&ݢ�����|x��Pf������5 ]Ei=GU��Ȗ(�Sϯ.�a�/p�����~ۃ\�{�T,���#�NUT�Y��B�m���e�����np��f�㭔G��3~��v �WߎR�Kw�C��P�,�}4$N���HQ��C��_��-��}�ఉ�FRʠ���y��&)b�y��)(�7D`�(pO�/�Z�w��U<9������@j�Y��M�P����K��eᚻ��t,����~�;P�����bl�l��fwP�B/���R��D�H7�˦�����P���Wev�׉X�h+T�Г�����
����j~���ԙ�f+���Q�f��ް�;g��d��tGܴ��|�y�6�{���z[���`��/+XQ���y������ߟ�eJ6�����A�x{ʹ�#�!/vC.�e�I�{����O�,c}T`_=�7'ȿ����u��>Ir��g���Ymc��j�� ��E�_�z�Rjꦎ�i�����'I�~s4�##��E] ��97Qb5�@�^�g��=�3���т�j���k{��oz�]1�7&�fF�H��� Ah�m)�E��m�^�
������S��z�jIZ&��ˊH�N��%����Ks��Eğح)�Gʙ͆ҴG1�W��T!:݉yЦ�Δ�/��x�S�S�x����^��o���Zvm�P薋����"Š����������qT��uR��>t��o��0CC:/4���@�G|iL��1}��@���h���×��gс��y�ѣ���ˌBT7x�`���p뾆¥y��Rpk�b��A�����_��d���k5M�d�^�����h��P!C��kn�߁x������񶖺����x���p_�Du~�c���	~Yn@�\�6bS�Q��)3H�֭�J�ܚ�|!�$ث�l+�k�N'9��7c��@=��X���1�߳~ޭ) >��h8	���!f:��X��A��%�l�˸B�B��*�F��綅��[35'a�3��b��͜��mb�b5��NOG���ʺd	i+G��Z1|�Kj ���`C�v?8ބ�Sڻ�
��:ͼ��;��-.X��=��s"�M_ ̪>��{���*��Iضѽt>f�(j���a�5T�.��O ��z�.D�B��{a�6������=����p`�Z�:��#�[�Ɲ�Ofo�!��U�t!Ĝ�`�oŁEYγ+V�B����(�ѴZ��o�9�Jdݹ���5�f-��NHL)��!M�$S��򿿗�A����둖y����'Z�ѭ���q/6�E|�hFk�S9Wb�u�� #��s���&	��/"�i��[9�v���5�����"�!!��&IPOq��ȇE/̝���O���Z��Ք�[{�ޣٓ�͹S�3���]Y�S��M�l�IPT����Z�!���M+��Ε��s\}�2�����հ��U8��ϿQ��B½���A��u�۩��O�^��5fw��Ƭ��%6$�\;�8�
��Q'�!x_ıza��g;q�=�6<e�k����
'�+�γ{�9�Ek�g"
�0ג���\���gr��94q�<Os[ܒ����W�c�[���Ǝ���9ݎ���-lr��a.4OƉ ����>r
��y>� H^9�԰�,O�5n�0�k�[iOl��,H��A�D)B�/ܠ�����|���Ve�Π����Q0wsDD$A�qѹ�B�J�jQb�q"�"�Q�F��&1ƅ�p��c|z�=tO�Q��(�H��}D)��^+�>wڨ����В������­-E��=D��҆��C�&_�a^1m����efV����<6��+��Ą[doY,kojD�!��g���/�j��n �a)=���n,
��#_{��(���-=���1L���dB� 8��2�TB�->���`��bH#��Ȧ~�JջT���hF��`',w�_���k=X��J�$�OG��L�y������[�9��~!˅t�	�<ֺ���_��5�#�C���ÿI>�InY�% VP���ٜ���Irn�g��2`o=[Q�Ң{9Kh������Z?���U��U0�Dx�K��~�f� ݨ�H����Z���=�������,>>�����?��p!�[�Y�������7vo'��	�+�����F'-EО`����EI���y�U�pP��F�tG����͚�a;!�:~����P/Bo�ܴ������ae][��k�w]���g�jO5�ϒt	H�&��B���%�d��*���E�3�$6 r���H���;���G��r�ol���qb�h^T���O�3~)�y��^�m��F��G�C��S }���D:O�3yu�oؖ�!(��cc��0�,��rí^D9��;<�>�n���88p�_��B�݀��"��r�}�x�:23�=4��zƨ ���j��ɒg������@�A�1�)m���4{�e�����W�]��D3��j瓬*��������x��#jbF�VΪ[����#tXJ�2lC�[$���#�=�{n8����l���[R�-�|JQE薼��\�����/v�&�=lal�V�m�D��q�UDݾ����(�O;ȴ6\���)\�yA�T��v��@����?���^u�������\U�h��[��u)F�{fR��šb�k���T i�+��V��=	8�|{4):��8r O�%�<�E�L��US�B�1�".�����`��Ԗ�-�o���j}�J�߆���\��"�uV�� le�09ǯ����n�ض���(���e�����tFРӱ;]�(��&�YgA噤�$���Ω�"�VFQ23>�f�D�!w�k��S���F�PL�`} �LwIqP`Rc}�C�x�uaR'�XY� �y�	u�?I!��$�VOl[P�������,�p.�1nc%+��2-�>(�29v{�� c�PlE�MKj�ܠ0�x^O<~��v'�~$E��T�8#|���$���E�_-_����0�xa=��&�\b�-z�l��i�׎�nh�#Xb���` ����|N��v��	_��8a�JkuP���r�.!4�9��q��F�� 6zr�8+�΄���.��]ɔ��̞��go	�C��A
�p��O�U*�dk��nU������@1��N�K�-ҮI &,>���j�D7m�Gh�B�7BYMjEx:��M�&l�~�B�P_�m�Z���7ܟ���(�]��D�(������#^{ L��!��.L��F�X��%�Bxbս0$�o��t�p淆��y�<��=�Bx�s$���YWd�����t�˯CE�����`Dh�P��H�A��\�16��NAX�+���xR�XG|M��[�������d�� e���b��e�P��Ksͥ�]�yg��Z-�o�ܭX=d>|Y��m���9�w���1�����i uݾ�Cs�bSѲ�a�Ij���q_��B-z~2�Ds��a��-+�U�M(�q��\e�Z_�����g���-Z��z�j��ƪ�3#Wf
����4"�8��i�������� ��0�
��,�%0g�P?.���7���b U�r�7��y�dR��7e^2�
�|N[��M肉�Pv��m��?���w���A�Ϡ��	�nC����~�A��
��?n<\u����0=���y}�]��)Xc���y�Z?7���b-f�����2RJ=�"ř��S��ئ�Aͽ�;R�;
#��{�ut�H�`�4m;��Dq�r9�	��Q����$i��y�k�ō'z�6x�DN�N�+:v��Wl��I�[�L7�6N�9���+j��"�Q���m`	 �"<X� ��T�w2��C��+�*E3�J	֣7h��j��<��t�HYg�\{K�G�w=�	���JӿK�F��N!�B�/�����Kl�����ǿ�N/��������񖲝�q��MN�`�Z0��/��A��2eoT��Z�����@l����e �nY���2ޏ����\���!�õ�Hu���2m����՚��UV_�Gf��ћ'5��x)��(C{ף�jlAē@ ��Dm�nz��iml�H����^�����t$�|���{��N�������Kb}c��$�Uk�������������ڰf��=��7�p����M+t�#Ǵ0bW�T���";����ٓ�����W�ÿU�[�-@�4	��5�R}�$r�b�_��A��4>sa�{<���x1C����)ݾ��Ja���Me��X�11�aod�D��C*�k��K�~ц��p�`�,���މ�F���p�ҩJCXi��q�s.�5�)M��S���^�����pesP^�wQi���T�X�|]��-�C��� �_�I���%�M�p��
f�ݙ�\0H��t��t�0��G��(�TC�[G�ܕ��&���Z�-��'显t�Q\i1a��S�����3�Yy� �y�(;op�7�t?TaӼ1Lݗ��|f��ye���I
��߉�r�%���i3.ɷ�.2�xa�k1�>�=�(^2�SMHq�.��`�B��]cBL$W''ej��jrF�����a��9�$ةO�����²3��r��\5H�e�5�dY��2S�I�>�oq��r��b���N��������x��=�d�b��b���I�YD@>���"����K�����mn(�hwp���ek�b�^Oo����EA���� |a�e�uZ\�D��R��F��w#n�U��u3s��A��7
�����ӓ:���������}���E�dc��+��PK{��z���q#����]�4�wUZ���Jf�r�Z<�Ձ�9�@��	����x3��e-X�I:�W�Z����uKO!���0*�^���l�R3 ��``oX2�� r�!�o��gR���<�j�"x1PM�}e8:�,vj��e����ַ���7	�6TT	��Y�°(Ѝ��"N��5;��X>a$��ͦ�Զ\���>�x='�.��n���R�`i^7G�)�Ǩ..�^��$�Qxf��k�����hWjv�pWqJ��1� r�Ԃ�'M����ɔ���]�tP��>#�{m�Î�Tw��:c�RR�n���>�ԡ�� Q�f���n0��˦�_�H���d����h���;�}�;���³� ËW�"!z�"��' ,vʈH%���l�cI���[��9�)-�Y$v��u4x�wE+����f"���͘k�u[I�16f���d|#�t͈�%��%bX����y6��OH�{����^eJ�V�V�IQ2���Q�9�����"���W�U����A%�sHа4�aenw �����9���ݿ�h/����~N�~HnC�j4Ӥ]�� 3q�byH�7�w>X-e�bn�bЍ��,5��k����;���\k�ĝG#UKa=�k�S꽹!��wl���0a�^m�aL�F2��-�O�-U8�\LN�#э՗o�Wx'�ċ �����l��%z�z4�2Ky t��gZ��n���'uBo���# �/"$0��Z�"v��h7U�#�?P�ސPj�T�@�5
i�Y})�iN�^'l����Y��u��/n�듯@����WpZ�PD]��M�$3��J��?�R(lj7͋���|+�pxt�
$�q��2"�2l��jAZ�I��k�@X|��E����ә��!�{��l���S~6�5ʬW	�BS�~�f������3��?c�y�������J����X���"�^�D~�����ރ*9k�ؓ�(_wqx�����:�IȒq��6�$�&Oez������r����I��٦G�zQr�H�ѿ���jTF��b^�K�]�7�L#��Ψ��Wc�a�N�fq��U�F�^�"��m�y��eH��}{]��"{�t�����׎n�`g�{͡����5�x�rj��chud��p��u��=�WK���[s��hfT��Yg�2+��B{�������x"�	��>��* �H�qm�F��02����j�m2�f>oGIc3Q��=򄂈�R��F�{��wr�F�׭������'�5� �M9��m(���&QF���x&^��H: ��}*�Fg8>���}�����y�x[(������^��b���7���� �[�_s$����]��j1)%� �9�+Ź�۾,��P�$���E��"JMX��z�}�k9H?)�e��d�B;k���HЕҩ���T2��b�=�0ͅC}��P��5�y�Y�u��d`���9�U������wT �w(}��� ���r1�9bo�YO�$:���5�>�: i�&r��Q�X�h�����	��g�p3Ƶ41�௩d�^��������'�&O�f�nX��~׺�4/��I���{�/
l�K	(M<=(�F�N���=9��v�Z6[��_��4Is{80����)�01��x܀��sA"�P��L�M�C�N-t1�����u���\n�M�W�Z6��t�_t�A�w<σ�!q�<���U'������G����7h�z;�	ыW�^��js������G��v��� �"wz`��'�P� t�8/zJ!Js,.��¥7D?1}���[e�#�K8Z"����#�[Q��(^���qQb}�5��9d5+�3��f��0hE������T�����a��mF���^g�{���_�.x_�̵��)S��].+%�����x��l����[4W�'��'���
h��նk�;�����{���2[�%�@��V�P79�{�_a��V�S�߱�!�#����Ձ��_�kK��9��9��D�6�=,@�n���	0�S_�2��
D1�}YЯy;��Zw��Y�1��u�*�.p�o�BL�e;YN���P�Y4�Aie���'ˉh�Ֆ�8e�(mdz��C����Y���t��(�����}@1с2�?����şK�%%�� �o��Jp��YI�Ò��u,� ��������7R�p�5�o=7��8?rR�)V��w�p�{�*`)��=֚Ȯ��΅Jد�z�Qx��.�gm��2�t��^%�v>�3~��2[;B�^�:�7_�����Mi�=,�<8�2�w#@��L5 �����IU�<��	�쪮��֧�ko����nc�O�ұ��v*�B�k��
�����7SnM�d�4�?�p۸<J.0}�*��R�@�M�����;��_�V��Pa&��>�/lQ�2IX�Ihߚ3ƃDSH*y��J����.,���hL���WG�=B������K��?�0j����W3YQ+���wa���`$��|�'<�AK�H��6p�2��3�v����]W��9zf}O�O~�/#+��SL*8�J�AE�PS_<I8�@��</����L?�g>�6�4�uKH~��Zl4��%GGN ���@k΍9��P���q�l�fi��鞃S��=}3廲R��F���zS��^�q�g�,�����e��+H`r~�Y7��B����`�\�8^��}�6�_v�<����"E8R��g�6(��0G�c'��:N����K)��"
��gd���V��wf�la����Y�"ǧ7���9M���f����	�Ty$?j>&I(V�Y�t�oEc��4�E�f��4>!2VKR,�ۄj$=r�ߐs&>pr*��,�UE���u3��ܱ������`2�S��ƽ�c5_&��	�D%٪W��ٺR�FB���5A]���FҧDGg��P������U��f�6�ck�����F�ڍ75����5��f$i�W�W�����Y����p���~�88����L��p��+��^�̳�I�2�}E�O3��~�|�JgUo��z+�/��E�ʩ C����7�����^�ӳ���_"�S64\�!�|W���5��E0��rr��	j���s��䉿Ɛ�h͖�;�B9�ã��_���J�Kz��
��:�N��s��+�H���ǝ԰~�7��ґ��3���]$ |�F-G,������fmM?{R�͑���T�1^��Ԕ�=�e��!Q���&�H����(n���u�s�iN5��+]�m<�e-#$�	���_tj/q�Ʉ���	s6�6�?�|�R'�M�����3��P�g����b�5Wi}�O^��:�����t��d�m�&L��2A�z�^?�Y�Vō y+zߜs)`���=��n�Er�{v��J���=E���s���{-sc&�Lo�֫'��Mk|S��[�Z(\����bqz���7@�r�%U��YBDͺ�Zk-�F1-5P�>�6
ԕ4�	���|˟$!O|	�Lz�H�v:<--J�8�#)�|����h�S�	W�J �ڻ��a*k/���G�5q�!�.�1�(F��K�ݼ\o+�7��1uf�w�,��G��YtO��]�-���/Z��=߁n��$K���ޕ4_���ɴI���X�ۄWɍ/�2p��~.�H�m7�{�V���s���x&.
p��H�<B���� {-�X�1�~��O�7��R/�}Y���iT�(��%���'h�qms '��b�P�T�h4�}I���7��|���R�#)��yWpK43���ﲟe��b6��8�(`N��z�YX���T�F!�O��je�f!!���:�� ��*����+Kأ�Yt�n��,�OZy��(�����z'�T3S,@��u8���dȹ�]��q'��X;o���˫�
,���̸A�v��뫢A_��w���r��*+�[W1�z��Q���[@I�83Mh=Ä;���v�4����وj*�U?g����r�������BQ��(���PJ�.�A��a��S�)���۹�t�,97�)S|�6(�(s��>f���DJ�0�r@=0���%���L�����5�΍���ٕV�|o89��3��ϘAU��(J�z&��i+kJ���k�� ������a�ЌznN� ��H���Q���Y*��( ���x8�p�f8�9Icx�?-ӒϟPKO�ޕ�R����D�*���ּC��$Ӽ)f����'�%6�M��İ�R��US�*��B`��7��JS��}�yl�5��zҜ��}=km{/[Qi?�s��Ɉ6��[1��S����X� ����K ���OSʞ 3�MM_'撒��^���\U ��$ĬCr�ƀG�Lv
�y���D�����r�.�l�M�^��3�"�GbN��mz,�k%@k� 	���l��� b̹�$��$�2�����a1��ݔT��A[�Ff�K�GAvlje�`��xΪP��lP�mT_@ι�j�N�&���@��D:��{�����qɩ��֦^��u�-��%�t�����r���'�~�f��+��\�y�s\.^�X�ݟ�f�]8Y�¦�3��W��q�.w6OM&��n��n�?x�K�� 0�2s
5$(����}�X��n��w���񓁖Yjͭ)��ݭD��F�1sm�R��3	���A_�Ώ?��<���>��<��3L��w�Ʈ�\�~�q�Ь0E�~�֡�`(�!�C�ϧ:��b#@��#;�����Z���Xt퓧�w/a5u���:�t��-���z�}��P�:≒+4LW�!�ؔ��r���\�ؼ�y�Ё���U�Y�����].p�p[�3�n��.�J��zq����L��U���!�9QNt�t�'+�-BPY�gT)� �y����JE�c�&���jJ��	����.˔�<X��uw���� �K���r�KS�cA�W�����t������W�nnʀ������V7��y�)͘��^��t�~���+6;��� ��@2�)2}���ˑf[V��P�\:�7#o���Zq�{u�����Ig�	I�:��h�̮�j�\���(��f��}��u�����fJ
�Gx�#_mh��H1O�
ՙ�_M�X�:�CLJ+��K>�+�*+���s�U$�C��YY����g�܃=\ |��d���q�0U�'��IPg�&����|��Z�U�k��"�u� � C�g��u��I�7_�=�$?��C�$�>��J@��ǽ?�4��cszگ�Si���<q�����L�è�&L<��DjT�����/��f���
=�� �H��w7����tQS��a;��U-N�-�$g*�]�3���I�ɵ��{��յ޴�|�2�R0D���HĲ��\�O�%�W�~��X�oȨ����%�ᇒ��X"چ�������N�Y�;�w�Ϡ��P�>- ױ�;𞌤Qh�dX�Y1q���Wg��'ۍ�b��c���������*m�6C�Bo潮U�:AJ���0S��L��7�l�����6>�j�Dt������yN2wC�@h�"ޕ�� r�O��:- �>�ݽ��b�zx�̓�)��]x0[������:���]v�=S[�"7���ʏ
&E��ޮY
��/H!��
�������g~��B������q��%.X�� ��t2X�����p����1-z�lg����\�>ώ�+e��p����z�x�����vvsu5�h�1c�  c]�wc�;{
�^s�KY<UH�>t��O�K��-!��l��5'����'�y8@�EA�~f�6���$fz\����
��^:��y������e�$�[�1P7�J�橤�H/sT d�\�:u�jO�o�����fQ؂����`}�jȽO�b)E�܀J]=3~��ʺ�c�J|{��;
�Y0�!f�����ŵ�.{<�ԦߦtD����n�{�,?�h�P{����R�T�����E��#�K�>�Q�:�cA��������8L���+��}�_�ڐ�)D`N>�ͣ��v̀yA���~�	�gŻY���
�O&]�_��p�_X�q���&���ܞh����yd��X$ᆌ���o}�I��J(Q���q	|���GZ.��)��ߌ��f�~��m�>�=��:����둁T��ڀL�]]�GBO4O����#�z��.�^o$��m��7CtЯ��)�lw�ù�	c`�o�/�2��9s��X�
��GJ��A���/Z���i�Ӝ��� �����~K?����o��I�]m�O�Aa���7^.���v�k�li=�m��{Wzq����`��ݰz���H�:�Q�K�c ��M�UO13?`Xm��V�)9���+�V��F��X����D���
�ߜ�$8z��R���AT2�l���9h��ڈ����sGޙd/�5z��<��voG�-jB�\�^�I^��KL �"d��kЫ��>J��6 �rGl�����;��:��r��-�y�h�[=�DQ�ꆄ��0��s��bQ��:78R��d�#a�UϪu����<�<�4N<�/�1
��e�������n�Դ^���}���y�l���K���.�,�l8�"��e����X��R�_rY�9�޲ �GK�\�s����LI�ɃO����r���ۊiY�Tg8ܷ>�u*q�ϐP�P&����H���KfΡ[=�2V�/���-�Y�N��_�&��~]�j�m�E����O"Xu��I� ��%��&xzlM��;=�����L�j����->��8��?��XO�	�~��E�j[�,� m�����6p�sg7��(}��Y�o*��Ю=tJ�|�D/��4#���d���坧��m����%>_RƼ�PNe��58�K@M�/�©��
�� �H ��D��}�.��a���Z��I0L&��-�p���o�p���䈍��aܓ��7���{�ua����]	j��v9��PX�����e����t︚OGH� z��F��|��8���k���=ΰ@HMY_�6�W�
҉į�6�Pln�潧$�K�$�<�i�pŨ��2w�r���~W[q#_��1si�.�`�Z�71�pkJ���?X�L�-AS�e*|��/$\�2�P�X�T�������i�͝ު؈�b���?��В���JQ��3�qP~������њ�σ5Й ��(��G|D�	S�5�3/[����{ГJ�c��:hi*��֓X��Zv_o��.`�P�Y#�}��J�f��"��L�1{�	Ng�u~}��2�OM���;�<�`?��喂������]����1U� >FF���R��#j;4��~9��đ�����ڷs}_6YJ_�{�7H�pCC0�c.n4k���Q���Cf	 `qL �V�cVU�_?� ����'�kD"<�K)�ϦJL����P��Ⱥ��m<5e����e�?{��%��!}G����F������K��= k��*TM?xv,�a�S2��hؚH��������!� ��ZY�<d����#�Row���4�08�!_�m�`���*�J��0�v� Y������8����P5ז�S4��F��jb&ͲC��^��jE�S��G����ى�["ɾ&��٨_�sPW>�a�R�B�M]��
��<�eX�ney^����%�����f!ɝP	r`��Y����d�˔���g��a���U|�\�Z����T��Gc����I�"��G��r��W�!�3�lۜ?�����7��U���i,�"h}��P��3v��W��A:���v��	�^��3KM�
���Z�+��i"L�lrV�7�,�����&��/����fm<=b]+���;;R�����4I�U�]�F�6�r?Zԥ̯�6�ff<��I����3=�רuE:��W-F�y���!2L�������E���� ��ckҬ=�EJ-X����O����a(	���rp��ֆ�r,ѻ�/�	������>��xX���r&��RS�?��9�غE��S:P�+�D��k�ȣ�X���RpG������	�g�	�μ�ء�#֢ �wl~��"��)�&��
*��{��s��L��i��H-z�z�C�=����]�JGVݶtX�J<�lR]V۠s��;|uؽx��M{�T��G5%�2kxz��a��KD���6����*�Q��A�(G�g�Ќ�]�r�U{S��2�)��C˳C����J�����)�,!�5�]�3�ĲE���[eI�AR��/
U;/��lO�>���N�'cE�K��&�=q%S�Bc4��XN��/���N��0��s6s�!��:��OS���ڃ�\��U��W��O K���&L���2$���pC(��^�5�Bn�5��\2���Ea��C%�r+]@��ʾ��D���-�n{��Y���|�5�%�����@ȴ񠤤J	�p�?��k�_��e�ܜ�W��=i�]���},�Fc#�,H�L+9 ��%��rL9�&�囑�r^�$��X�?[F���ȧ�+�� XŮ-ɉ,���rN��rV�,����l��I�@n�ҳ_(=��]����2�a�m9�W�Z߾eW���+�	��-�f�n�T���`6L��EH��*��p��_gD�uF���Tه6}�q��N�ZC��Ok�i��1<bB�~٘L�l��gX�P����
R5Qѩe���B�7�7ۚݞ�]�3���8E�l	)�� v6c:��ON�kacn]@ME�%SE;����))JX�x,P������N���^DxS}#���H��5��ˋ�{�B������3ؓ9S�)X��~f��~ ��.�2�RLo��Ya�w��n�Yt����� ,��'@)��u�`;�����cۥEs+k[�@����#�k��̇�\�n V�LY��R@=omtWz�P*�����C��!~p3�M����C$,���-����a�	���=���k�8(j���+SJ�d���I��uM/c���vC�S�`�6�E��$2� ����{}ڳ/�͈���H�q���4]|t2�筗�%k���ᄗ3�TB���!�Wʴ"qҭ蚴󆤷�RCa�"�]~����@^p����P�Lgr���Ʋ~������H�;y!��NKpM>�b��H�[� ;���E^�P1/S6�w$�Uq�/���2d��ظ]�વ�K't���:	��`���<Ȗ׊����8�2���lN�;�#9�}L<OrăDC8K硖R�J��9�ǄR��)��*C*M��f�{+uN��P,]�'��?8�Ƚ5QU�oE���旚S�E��^3jC�ț���L&��g��;�ʱ	�ͦs����g߽�-��%#��v�l�k8��Ջ�+��D�_ő�%�Q��b�=S���7��JG���BeOI����/�`������!�H��\<*���[�o��{���΄�G+��ѝ˼!��0ڽb��&�(Ж,Q�*�I�*5v������X�=~p���� ��unFs��˅Yb�e�fCgP Ts!F�P��:�s�kg�1ҧ{���Z�;l��x����!�E�a�]��C������O�K��A�&^f~5( kG֥C���t�R�˕Y� ��\�'���܊T�te�,�[B�j�ro@A�H���.�cȥ��z|3�wS�R�`ywi"�D��:�J��ʓ�f���0��������_׫oU��Ӯ�y$Yz���������Y����d���dl��w߿�U ��BwC�Z�-��
��}<7�U}%|�~���^�����M�3L����qc�L�r��l�!g�	��3!��v����β��<;�m��+4�@��ɥX�C���[.��AJ�4����mp����):�p�w�QP#r,V����s�H����O�nH�J�+${���ja��A1�I��f�)�wb>#���0b�<u����v	y��#�a�ic�n�,dWD��������1	�Z�i)	4u�DEla>����X`��6QNr3Aw�1��i�7!poFO�5���h����P�f��*8)ZN�f���¸-E,ޗǳr�M��Ĺ�U5��0HD�K:_�b�������"P����
���7��Z��8 �e����M���(w~�tm��vv��6��t�ȧ]�ib�K��p�

ͪ�߆�]q}E-���Gmq�S�>;#TA{A�R�¥�3�J�	�*?Y�f���5�r���+Fi�k�7Lo�gگS���,N�+��/�6쮶��v�V� �v1d s!���8D������L����E�М�֖jm�2���>��C\ڶ�tƯ��\;r��NL�%�L����}8�n�a��s��Wx�������T�+�PPcR���J��-�!�d�[��]�0	�]T�\{��MH�gO^�(y�D��ю:��.�%4��O��8|��y���fT?���4�@8�Ba�c[i1�o�A��Z�T�2�����M>dڸw1k�+
��E� ��ڙ����D"���[F#��%P���������+���fs*Z�
e�Z
^�з@]Jʌ�Zt�W�c�:�r7(����ylq��,��t�F��8J��NИ�'P��0/��Ҍ�;�"aq�q�==˴�"a��Q����V�#f�����-�f�A~��%ε� �ڏ�cDj�l��<��f�]���	Z�q]O�5�*��	zc>i�ئ&��[��F;��lb�G��J,U�g����A��9�qL���J	n0٤n�Ϧ��;��=G���:A�'��|�:c�#7��Df ��~�Ffa
-<˱*�&�5ݸJ�3ā��%�L�4*ZJb�n�|�X�z|�QFM+'��F���7�ʅ�L2�����=����~~�϶�9�#o��A	����@������Ȗ�9m����Od^�'�ٷp�`U�$��95B"1�7�Z�`E��hy�cG�(�H�R!�R�/�<L`rw��eٔb���ú/P} j�ft��4��0^�CK���̴�S	tEl9.��¨.I݉Qd�p��+֦N<o[g���*�z�>����t�~=��<~M�Px�ax
�Kv������+}��o�h���C�J�S�b�h#�Q���+��C��Y��Ĵ��8:�H�{�TzzV�ѕ1�NBh�ފ@��7�.�=gwA�L�FUv[�%�tu�"j�T�];*X0S-�l~�j#�"�g��eK�������uUGу!n�ª����)�k�e�H#����������[C�S���,�w��L�J��ۖ!rf���T��{�u��s9��	�3$m�1�vP����� I�;m���juf0��D��a~�d.Ց`�Z̺��hU�`��G����26WƦw}�W��n�ƃi��`_4);�������Bb �|���#A����������Ή�>�T�Tg��R�i�7�D4��eN�.� S*)=����F��O������ո،}�FF�n�I���.4���U]ۉ<;\��)c,�s�ؽ�dP0xQp���Um�I5
�&�Y`���G~��ךG��D���o9�#���-Q����\Кf]��B�j-�sr��i⸁�i}0�M�վӊ�9��&��;�EZ��� ��#c����?~�$�)Rה�F ����,�;���wĳ~S��6޷��M��j$un٣��u�fw���QnD��j�b ��?CF�L��+R��*�^\`�`�ՇP�l]�����U*������9-�t4�#g�
)-�eCc�d�tl��J��U^�sv{
�����K@�1��zh������}�+1��=]��ӊ_?Û.��bp��C\�V�0������a��}B�e
c��iL���r>����+��VR��q�X��F#��#��c}�7��=��u���G%��b�k��ӭ���h�>.u� �����@��M�\�	�6b0�H�O�e�x���8 ���<~O�s(����$������"�1����[�6�u$��*DW
��z 3N*􊏏-��@�x$��Øu:�@����x��n2�Fӻ�����a1n��e���Y�9�&��
0��%��ԋ�}��9(�+\}��XcI�B�2��V��B�u9���
�
�qؚ)46����=A���`��d ���<�UG��79�'~�fa� �Њ���+cg8ڢV�����@zԳ���}&Қ+�X� �є#i����m��;⑔��wX��M�D�;���*Ƭ��A�D��R�Z%���D�t&6���8���=��)ϢL�qN�����EߌY��[*J�~��,�>�hJF�͠���\6�byy_�t���k7�0��,v%���{�N�3џ#� ��ZE@b�,LŸ���~ҿ�AM�V��3���q��6�����d0�H�A�С��m^g8Eg<9��G=e�m7亘�\/ټ���z3ѝ���,Z&��\�fhcM�Q���٠@G]+tS��F
���:#�M|�y�pŢ��JF�����SwA�w�-BM��M��qd���W���s�(̑2n�kQ��Ͳ!Ʋp��%`9c�ٝ�DR��\7�f���;5������(�f@���8׀�-v�#�U�b��E�Y�a��'���Aa��:t�%R�. ;B����������ǋ�a|��3;Ҡź=�c	��C�z���6��l�=�_�,x�*�027�5��q��S�Z2����r�wm��;��^z��v�^-.d��s1�$Z7ߦd6���{b�_a>�jܸ[��C�k�}s�'�=_�J�g�
s��sJ�*j�"��Uk�*�$~�2��lAf�b�=�)�J/n�N?8��x����oI���cX@"��(t�|q�����l 6�|cI?�V�8��R�-:��FO�?��X
H${�Ln��šY���������5�%��}�k���9{5��}]L�&�hw@�u�xA !$G�� ��B��XO'��?��������;Y՝S��12caw0��lEv�A��i߈�7�
��Ϋ���ڿ�I�H�+�j<L��͵u�[s��W� ]3	�!��1rqjN����:�$l��v��>N�}�(��w=����w���zM�~��~�KT�q��s���x%��_ó=�g�)����LY��E������Iw!��:+^�(��ZB�Ց�ܐ_�ic��~d"G��v��3o��T�D��N~��]C��z�o�6!��d.�e�tR����q��Y�7����� �/4��v�V��W"�=��A:Eq^x�s*�i��t����~}���S]�j�VLzA<�?˂T��eC����-YW m^a?��ؕ�񻹫�е�dT������pX�8ԝ��.6�T�y��.A1iˎ�C���I1�4����t~�ד���I�f����)Ź(�Q��y���=��Ғ��
ͩ�Z.�Y�x����K3�H�KC�#�b�w�d�+�d/���H��
[�]?C� �b�,]�xР2�,��eF?yV�lKxv$�G����E��
��ȫ6�"��E��d�^�m�K�<�{��%�J'1�l���4�Q�#��U*M�>�K������?��|��
������5��>��="`�H��ֈ�Z�I��c|)q�>�Bp�H<�Q�wȐ#m�d��
@�ڴ��)?�i2i���`#�ˋ��$1�
=N����s�hGOk�A�0A�t� N�v��Q�Vю=��!�AYV�\�=�k��IKW��G��p?>8(���L�6M��c��7h��ge�\N �W����v�^b����Y�����ǎ�l���Fq*v.{���h<w�F���,nYȀ�W���>�TCùN!�*ڊq�2��2���^Z끍~@6o��@c�!r�9׳���lmXXt_�Sƨ�.�K`�"��si���b����-��_24d*�oeQ�$!���{W����E�z)����rGur
ś��!��&��ߞ��"Eu�\I`l�ݷ�V']����~)WIU	T��t�;��W��R�?%$�2��A���xWa����x�����0�o��G����Ά_:�7��[��1U���7`���Y�Q�)���[K�bh�d�q����,2�L�wjI<�Zc�)d��T}ťTR���r땆���,�Hb/w%䣸����5���^}X�O8��w�s�䯙��f�ÀaH}�>����c����6? �%Ss��&�7B�f��z�v���'�Ӹ=
>�P$��!'d�ܦ�XP�:|(��R�!�0���|�OcÍ�d3�%eb6��Сԕȥ�LCw��
��/���j��X��N�	��I�D�>��]s�to��&=�q��(%�\���+�
����`!���̃���9i��S�H����g����a�XOة�)!J%��������}��{ �wS��hfl:�Q�y�g��"��?$F�>�͊�G�a�e�^AO������! K��b���#�~�Ǳ9���v���s�̣�t3ce\/�GX\�	�5�\���:��eϮc��f�>Z�RC�dev��W\�X�	�q�.�H�oXd���bx�2
,�3RˬwP���mC���'��ԔʐA��O�H-���-}B �B��u:=�YuQCyl��Rf��p��N���9}���D<\\,b�F�V��&��H�"����?D@`�rKr�emx�&8���{�sh��ч����?��J�^"�m�	�I/jԳ�2��D���z��n�~���)�[�0
�
�]CD���%GpL'.�|��c��l]�L�~�H�/�cw(�BP����V:*���;o��WZys�����:b�1P}�6�w��qT_��G�avrX�զV��'Y��g1YoGF�L(S�SR�:Ѧ9Kȫ��!�Map��'U��=p�hA:G8j�LK"h��P�_Rbkk���MA��M�u5K컧�ky�@��ɾ7��D})�W٤`���lSA$e��|�.}�[�Ye�̾��� #~_4e'Z��'���A�TF6�!鋆�*��T��ڑS5��7�U?�2n"�0GZLq�Yg_��)Q�J���\n\�/R��V�J�*��y1e�i�C(i�����U`���ce	�����Tߓ@��~af�P55��ͩ�M;�v��Ol�b*��fu- ��:����%v�D�T���ᘶ��RP��s����<�Jl&c�$�¯���'�9 9f)�"��xW2.�H�����턶�� e��Ύ��#0W���׫vӭ�h2���?�l6~���m#�0�m�o�z.=[����A,��b����S��$`�&��P�(�fQu��z���m�xr�a�L�/�(M�Gg�O��K�$�Ba��6��9�f�6ݴ��y��N��t@'��|n�vB$EĿ�{Qa?d���YL��܆��:�_���F���;�4V�}gT�*���2J�3[ج�����h��#|�����+�Y�R���c��umR#G�<.+xH�)�+��X ,�j,Lљ�Roc$�b~�Sc� 2w&�������b�n��D�����>>te�?�<Q��#9���c��@P[yk��<�1�L9GD=�+zpɎ�Ao�)hZL��zE�n�9}�0X[lUv?�0���	"��k*ƫ��UW)Į�$xQx�\h�5;а��NP��cX܂ȣcg�G��h���5���_n2.=�:I�9&���@)⃞T�>�7,j���^16W��p3�!�n/�Mq�y4����uU���.WD0�A�Q��ނd(o��S�\�{�1�����WTS=�.H���݆��� �����p�{�Y��Z&�3�:���t/�<K3W{�
��a6©�����D1�&2��쳤�a8���3�>���ۏ>�)��1Q�ԏ�>�=�ԋ��j�л�<�d�[ �0vT���ʓ��o�~�����=��{�t�#����Υ�3B���?�f?���n�<�˝D����7��O9���c�5��}TrBg���X*Z6s�zg\�䰦�E�P1���O�¡AM%�h����J�Sѧ_�S��*Yӓ������*&Y2�ou�7�J�Ӻ���	"��3�����# �7����X����+�S�ؼ�,Fw[8�"D��X}R_cN���G�W�IZ���+�Y�4�|�D��f��O�g!�l�Թ����@���2%�Y�'�tA�Z���u��}9Cx�����¯!�Ac3���AHA6��Z�zm�,�X�g6@��޿G���u���ϲWׯ�!ֈ�W�Y��R�mHE
�;̭��迖�&c\�
F�
�r����������_���#{w��N��hJ�pѣ�k[���#�C��x]\n��T��a���_��w��g�X��1T��!0rzZ��bu�+��3�GMB4�����:��I<�9Ƞ�{ʃ©���H�BE��L+�FbGp�)z�`�PQ��8ޒ��lMH�R��Z� �\�ܞӵ���)W�o���� 2��;k�@���c�2���r�!2!Xw-���핌4ޟ�d�(��%w�� �S!��Ë�A9�_fy���F�K����h�R��8�"� �|�7'ϥ�����<`��٥'��1I�����AĆX�G8��E}�'&�&�z�����MD�v%�{����$u	��`�I$����SG�I3����-8��U��㮃�m]�B��:/ł�$�6���`�\����Ow��쩋V(��)#X,��x����;eͷ8���dzz����g��^ ��`^>�)g�5嚲��B@Au�a�r߰��]]��ʡ]��G[�2�������Z}��������H� �un��oUt�d�2c��^ߧi�;����2@���a9C�Y6��B�j��g�S3'墆��d/�Z1M������e�z�rE�M*��� ��>Tѥ��m�\�)�F$1,���ҽj�������d4�f�XI�ӱ�ɦf�
�+��X	�&7���_M(�O�4CQ�N��J�C���(��dLO��\�5�ݣf�(��K�o!�C����#��y���&�TO���&`���'i)�Z #�7�[�^��f� R�.`a�]<�X&�	`
���e�bg]���	N>�/)�'~V)}�co��Ѳ�*=�Je�����+���U��6��OF��;��.N��6��ڂ� lE,x;Ŗ�q��R6��!��y�jԹ��Ft�dx�c	l�TNU	�����[���G�w{6��Zc��v;ފUO�����"����+���5,��h�sj�'�n��i`w7\���8͵ڸ(��g� )bf�x(?#��
L��~!����Tٙg�V�[��CJ��u�!�7�`�a�����:W���������Q����ʰ�R�<A98nA4��a��_�M�-�7{�"i�fc��=_�){Ɩ��`
8PH˘��e�G
Y�W���q�����Ǵxs(���.�qL�IJ#�<���W�!�c��PR�|�X���C����e�ޢF��XH������D��=�ÊǴ�C�f9��c����^��\*�K�J�\�9�h�Z.�����L����� ^�ܾ*`�/�s�r���v賜�zi�	f��Z��
� oI�o��=v�
*+QU�Q@h�,�j]�moEJ��(�&����7�¬���/ťc��~�F�!�Q��PZ�s��T{�7���>v���x��5c�FU��t3��>HH�����ߐ@��8�,O�<؆��K3��y�pE�Xc_z3"����0]����&�a��sl��wvO�f�������:�V��l��Ucy������ٌ��jծa��Qu2}���Ęy��m��+�ZaXദM�>�2A���16���vP<S~'�5I~�و����ߐ���w\g;e�G�H��gC�D(�5������p9�W����)�;�;>���f�l��Fa!�b����p�_��I�O��z'sI��;���h�@����U�G����K�P�[��ˡl<,���R!�%B��^t��	�g-e���6�͟mk���s�����C)*��t�)�~�ť���-x~��WK�!����Bx(��'t��IS*3�7�H(�w��t�ug����S�#�-���In![��st�=���h���j��a����]�Q�3�/
�z���y=�ƅh�%����Jo^n�e���v�#	����;q'^O8g'�2����+P�����c����u����e1��>�����<-S��f��b�u�H�w��X=�s[$�\��y̠ȸ�0-V��땰O�	���!%�2���b��M0�#u��!ȪHq|&!�3��4�Ld�t*��N{py$;�_�(�綔<^^��X�$�c���-�ѽ7X���N�w��;˭�.�:.���o�\>�����=%1\s#i~�7�J�CR����SٹK��;�<��E3��E����ʘKp;�z���A�^�7�m0�w�w����ҦvE�:���	8�$�X��t~�-s@c8��*U���u��3�;��+]%cQ)�Ӫޠ���!+�;]�	���Ņ���+P8���%g�w*^��@!b�C��(�M�g��c������>��OG�Ҁ��1S�*���{��ЕrzRQ%��� .>`"�u\��0`6!�����õ.U�܄ER�]�l+�+3q!v�-j-e����Kjw�WU��x���3́{*,��f�w.p8�h$
?��(�K�Ď-�p0/Y�ʪR�����e����AX+?��\T����Tpyb�fz���b��
T��R�!>R��Y�;�2��1)� ����/�g�0�v���`���`C����r�9l��b���$�G����,�~��uA�	�a�_��0� ���w+�3�;mg�����1#�">���lX�'�Plp���"��V2A�O��*�t�����x�X�����J��z�j	�fB�b�:�٫�1�_.s�������j��a03ю�BV�VF�+0���-:�EUyͼI�h�K�B��O��d��RYmm3�\F�)P�L�m�}tg�R�/��¨��r��m���4LT:γWl�g��S��<�V���E��زϏ�X���Ėx)z~i��⳼M��BY�_HÐos�����ɬt�����T&��-rs��w$ ��ޒ��Z0xM���KξD�$������  �RZ ����Ü}&H���C��@Y�0��{�U�����И����=R�8��� ;t�x����<alǴe�$rP0W����ޱlB܁��bY�1�+��T�y^a�}ĭ�E��!�]uEG���`��d{f�1Hi��/�d.)�����NLAE����p.K���ey99����Z����`�������H��8���\jH3S���B#+�"Xgb�`��p��d7���i\�Y��K�kO�=�`PǶ������Y���Y����<���hK���@į�t���s�4�H��穈�{w?LpԵ�6�r��d�O1q}!d1e���sq$�'p	G�\��5:�6C9����^��o;u�9������y�,Ρ����Q,��EW��2.�eN栉�Qν��%Pw��e��%��ͤ�Ԩ\9�;(�����s�	�m��>	Af�2�ؑ�96��˺�\`r:~�d��jҞ���p~���P�Dس�h��i�e�!�X,R<�j ��Dm�p��(�l4�K	����ʫ)aK���WF��bPl�c���:�_�m;�� ���^�:�	��
�WR,�ӈ�$�����l	yx�4н�)�+LD����d[��|j�ȸ�p#�O�Ȃ"�7����<zRD[7oW�ˢ�� h�5M8�!D&;��'ž���lxU��OdS�ܷZ\�L�K��v���"˃�	㗴�v�mȣ����u�k'�N���ƬB�.2�3F�.�=Z�(ډ�dwɟ���ˁ}�F�0��{������9�;��8S=IZ��e��-D f0�}������3-�ĕ�J���W���J��at���`a�l�8ϛ�C�]f�� Q��>a� xhj���'����ll.����m�v��&GL��?;��K�%�闡9��t���|������.�����@�\?q˒خJ%p�����ϒݳq.��	���&��|(��;)�����~7D;�v	��?S#B�i!�R"d�<��nrί:��%���ae5Yf`�P*�<���.u��8ʓ��V���ٹg����|�'�F���*,	��ĵ���VS��� ��N�;ώ�+�W7�_�~�²Q��`�&0w˯R��[q;� ��z�ω��o����r���]>��������%b�su�G`Zޠ��.�|7��AY��@�m��iٔ��;k�4	��OVe��:�K6<�;���JwW%����
���[䊓+�_(ҡz?Z�i���tf��06�0��f�n�R)��@��{1Z����s
m`r��̩(��W���n�J��!����X��ζ�z	?�g�$!�\� ���[^��>O|�'�eBs����7�PC?�K�e5C%�/�~��Od2b�ꠌ���J�q��IH�_ �KL��i��:h�Q�G�R{�����-b����P��T��=��	}��A��]���e�S��>�L���N�D��}@%������]�#�&5�丹�c��gӯnXu1�u 1����q)APb�D@�bgTc�Ÿ�`*Z�a7���Ѕ�m���(5���q����X�����ID5�r6�n�E;ҀS�i:J�Ԣ�����$6�����k<����O(M�w�e6��,�A�TӀ��Є0@�F�l^��쌨F�8�lv���Vگ/ov�)�̀Uc�N_����e�y�Z(/pՉ�����'�&�TU�G���dn��uk��7���E�>*�_�w�[ڜ#�I�ϛ:s7��e���*�g#�R�}G �!:��?Ų葾�5;U2�X��I��3����qKE���:>`Śo�8��9ҥI�vy�X�W������/BW�D�F�>4��_������O��o�(1�U:���-���4v�9�wm^���'������R|�=-�8F��l#�l����A��H�ۀ���c��W@u`Zc���Fׅ
�Y�=�
�i�D�w����~��t������YsQ��yks�s2y�a��?��Fí?�y0��ky}�Wk��Ǚ�����e\��_���9t�+��Wx�n�(d�;��{h��$�Z@����@�Qo^]��/�"u��:ɴ�5>�rP�K�����ª�,V��}u��]�?�y$l=&V^�ŭ:��_\�o,2#�g><~,P�%p��W|�K�b3������Ђ�J���������	�3��IV����:��-@�y���ڐB�Q��Z�)�\S2C���1�*텓��g7�t'vXV����
/��-�X]��&)b?���
sLQ�3�U]�Q�h8�/~��Oss"�$bP6���{���6R��^n��k�qN P�g��Ubh}\X�F�D�0XH�VA���T�w��YÅ�0��L�=Y��gH?�e���AM��֙�H�ŪW"���F�!�9�㫲�����aЙ�uf�:!�B��� �[&B!�ԗk�R'�I�~�����3��fm��/�R�\����w5v�ȉI��I]��� R>�M��!�aG:�M��|\B���&��Vt0��B�XN���W,}�S��A��x�B(��&�D�w����	�F�I����w��tT�����ڤն?�SzL�&�����w@��r+�c��y��(��E�`bu�a^��� [~$�}�Q�`ƶ�����CQ�}��w�t��C�Ո��ö��&8���� ���G��_��6i2L+U�:�8�jP�DBE���4���\%���@��.k�&i�\94���ucuC��Ɓ_�k���;��h<�uF��Zt�9d�X�L	�� r�Л��P�o�`�2r����&����wG��
����y�CY!�I�sc����,9|rޟMB�aVR����zX��"��P�G���K/E6M���&�@��IoC�|P@'�Ho?��B��BP@21�!��Feď��(*� 
ww�4��}xq����Vjq�!��ǁ�4!����^����Y^��f�5����'�Ȫb��vyr��H�_Տ銢"�6����cS,�s��.Uri]�s��@ٱj�އ<C�#��3�^\@c�9�VS���&l���$�mp�3VX��1��a�k��ր�죺���&����DА\+>�|j�#{.i��;�0��`��gy/(W)� R�6	2h�=���Ph���5�o�_�n3���hh���J�t��x�c���N��K�����W:x��x����]ڹd�u��0�����'�C
?�dW�R�����]ƶ����=��խ*�W���9��=X��g�ne��Uj1� ����>���(�ݯ����fS#�#�F�&�Z	�z�$YQ�A��H}p���sK�%+�gf�M��"�d��,��(��+���8�:��%j�ӥ�K���_�Lyܘ�`�������
+h-�n� Rh��J/U�Wr��@�d.��Z����P���FvCu}L����<߾�t� �b����te��A+�9p���Gzi�O��\Ə� ����=z6�źu��a.n��'HÙ���W	r88���u�ZC�H���6"���E�/7�~bM����g(h��DƂ����\�^^{��=��V>{���t�6˲���32�eX����\ы�����<��7��93�e���򣏱Ǹt�v��9�P���@��@��t�_l�h�gD�l�킩�o��'r���~e���
z�-c������z~�����RU�3���l!T�t5�z���k��6-�2b%���J������g@�[Pؾ�r o*`&"]%V-�z3G�C�{k�x�5��<�[E5�K��*��t��)���h�����MI�I$H��vQ�ZķM~�}�fۅ�a�󂁣�*67��y�yn�%ߑ|��'�gy�/;�$����Bk�)���c����t�H��g��R1���x����c1 ����3��P��:d������àjf��$_�,���fr��ŵ�vT!t&4=8hψ�Ӛ��<�k�YZ�������f�������~l���?*k�@*�L�fਥ��,���a=�Qf˗Wh��(�1)�/��T����&��w*��J�<�Y)U<���H�D��]��29a�>���Z��Y6��Ȧɖ���&bE)I�8��T�F7O<T����2?2{Qc�^���%zƥV��jN� ����Z�[u���������6�H_�7�2'�C.|��&P���e-�5!"Cz�V���!7�ӛ~�y�� �7����Yz�\7�(�7C����L>��~�hg-��H8�v����M�
tF.��  K���$��g!_}�0�����ab��8�޾�`0���t�KtNE,���ɏ�@��(?נB�OE��0��C δ-���H�\�v���)�8e0)�]�nq����WƢY��] �*a.�z�1	=�;�x�UƗW���J�ʪ�k5R���g��ﲵNw5i�K����ޓ0nv'+�1u鯗���)H)���ľ��j�Ѕvb�\�Zz�5��5&n_5� K�k�%�uq��=�%��M ��_2��خ�,|�^�Y��g��>Ts�.��Zׂ����址2j��v���@��W�R��*��5\@g�2ކ�6W;���9|I�^ޜ�NZ�@Y��\(����v��N�&Z��L;:}Szfø�U��V�H_폣���1U�EHž����9;Z��1yWj��1:�MΕ�XM�*�iӅԳ!�������V�1-�̍ҵ�<�8�+a�A��^�T���w�^+��V���3��4,��dD(48� �4������X}Co�w��$�Y�t+<=z�?��>:|�%��"���~�(��G�[w:-�9��Z�q��1A���Z �q���=ޔ���Z.�ρ��V$�l}�|}�d�N����V"��ndj>�5	ZJ�v�k�a07Cj �780^���|B��=b*�A��-�L��F��:����H��'%ۓJ1S��v2Q��qW*��w�v����w�v��T8"�qJ��i�m[���i�U��bT�9 ��:Q\�96Z*=}�ꄴ;���19%��R,�##93��p�S��lJ�Cs3ߔA؍�����7R��Ʀ
(C��ؔԭ��UT�����}a�W3Q���.�/S���Z)u�׉����rk��w]�vn���u4��B
\k���INŐ9�$������*�~�8���aAM=��q"��$����� J��&ȵ͔+n<�)����l&�k�@�L*�	l�5.�:6�1�s?�2�=_��^3R9�z��CF?�����0?T�X1ld�F���<�>-����gJsv(�w�I�M��0�>Β�]��8Kc�� ��6{ݬ��Ŋ��r�*�e���le�%������3�g��ٍ�!dÓF�� z��X;݉�����dx�r�(+w��Jq�����1��J���Ћw���s>�6�]�&��:�H��jH�h*L)�\�8i�K|~���H� �o�j��6���.L_D1�\�-��/	~<��f@��-Ӵ���QϦ!�"��y�:!�zX8,|J77�:[�O�ԺT����<m� W"k�;Nn���?J"�')}����ມ��m��7�5o�>$�-����yP�b�	���V��3'K��o;>au��J��Ĳ���#��l�'hC���Rx7%v��mU�)/����T��˶�l���%�\9���8�087��e�{|��&���"#0+,�s���˰����wE��qȠ�R��EQ�<>���~�_�U�Ը�L�����QQL���Rm(�0��L�iy�~]��K[�BzbIX�*'+xT���V��KN��.w�E	!��?�[��������4��)���6�4o/Ͷ`��
*{��A=2�st�Ndxe䷗�h�B뺕1�Ul�' �-ڢe�47����rŲ�����0�76�S��^�J��
�eK�p�ա|S�����!6	v�7�p��K���v�|5.��ɦ�cf�b��JlA/�W�3�S�.�G�����q�ܪ>Wm�b�jF0K..Yh����h��!��*�"#�CxT�y%݅3[hZևx��h�M'6�� >�8�������� �R�U��A�x�F��ᡭo{����D��t��"�q��/3��(�O�zr��\~'(��V?fW�X��)'�t$ai2XDS
�Xt ���N���C���g.��g&e����!�cW����v:ѫY�y��	��:o(��f��q�pf\�s��fc��ɳ�h�}�������˖U�lPLK2�4Nߙ=�S�����t�><�2�$ +��' �0s��D��,u[��g߳�-{q<�DW$)t�q_<xXg�^�S��:T:����Y�$+�t���МP�k�-��\��eY��V��'���J_�� ��_����S�����*#���[�6慳�l.�z���\�2�}-m4[�@Ֆ3��2�t�ǳ8�vC��+��#5���6&%۳� oKq
,bC��7�b�-:)$��G)qsZ���+�vX���?3뜲W'��=,�T�3}��dq�c޵Re�1LtX�rԓ!f��A~L
I�S4����*�E���	��ܷ���e���֔���3?���[�B]����.��F�Mh��1��
����������>y�o��t�p�2��������T�6C)��W=��ys��y��R������!k'��L( f��uv�Lp�>M�2彍�F�m�.�b-{4���}j��~^q�Oڤ�Q{�=�?�����{�L6<�̭�LϹ���^�,���f�=��&��x�� �����|�{�EƕYU���^�ְ�r(��O�f�2�D�L�ПUU_> �*���ռ��MN��ז����,PWJ�ƗF-�m��a�/���S�2�<�ɿ�W���5��{����1�u����<�]c��.V�x�CL�r�$���,�0��yK�N�GbQ�*�2;;����)*6���?��\�
v��B q �ZK3vo��m{�p|Q�;n��u���5�CF�\�3q�6�$_.�?}ؕB7�cy�7��)�(�sH"*�хM<���'O[e��r.[�>�i|�c�|�/�[<�Pt����?J��M�.�x���X���m�}M����"�:n��qե����&�tJA'����Y]���d��-�RZ� ;|���{����>�ET �ݾ�mZss���^�R%t��<�R8 	�[�n�3�S�@,��U���:��MhԸn��8]�<���9��A�<f�xt�=�.Y?�0b�)�p�Ow�K	�p\�ޙ,�`�Y+��  {N�H.���c:t�)��ܾST4��q�h��R�9"�{�N�����sKѺ ��.w�@���E�:�f���}z����j��Z.E	O�}��("$��B��2�G��b�����'>�oC��l���9˶��"��]eaKz�}@M�Ԝ����X���j\W`�3�$x����Tw��"�%&@w�I�{D��o��C�M cL�4�����Y*J�i�=�$�:k79D�L����6��c��?���9��$��!��o���wi��Ց�P8�2'Fy�x�Vր�Z�;F��|��	�n�����M����<�i�qVwSn&H����2㷘��n���G��{i��L�sh��)��:I�6��q(^�D�.g�C�(5��e�*�&_j���jXtjH+4r�}�0� �W�:(β�ܲ]q����^��l�i�?!���`
A�đDw��>[����b�h4�3�A�!#ޮ����%�챟�REj �=�i50(6����8��'d��DC�tr�p�E
 N@���5q2c�.z  �:���܏���������{hT4�<����Ɣt���$|'l	�Z&-�+�>�-���.�^�l���̿Oo<^C�U��D�U_�C�zL�PR4_�w�`	�=)�H�k�O,�o��z���sZ:@��o����pe�ah���&@��"��nCe��?��<����������������vkb����aC-f(�\lC��H	��vzg���j��m�?��ͯ��k���wd�3&ԻT)��S�Ĵ.�x��X����k�X#s����Ⳙ�艭vd���qlSԌ`^(�ywr&�T�O0�����o߫[ɩ�p�w�|x�O��uG�<:�j��L�Wgo�h�����u2��6�VIZk���0��n=A�rpT��+��QE��j��σj}�˷t"�8�o䂘"Ғq=S�],2�tj!��h�����c�v�/�oH�����.�SHA�� p�7Vm1#�\��Р��(�#P>(v��[��;S[MY��	LI8�܉mlu7>��i��]ٮD\>��X�V��2�5�م�Q�M%W?�'	�\!X�uM
�x}"�q�A��﷠˱����P��gaҐ�e��W��"�i�->,x�8k֨6���ho���}ip��K�
t5��֦�۷�����9�IfEeX��6D+�5�nN)��*��,:���P	��Z�7����	�.z�;\�Vr����5}
�0KBov��e��dO`�U��+$��-�W\l��)zj/6,�ya�ͅ3�m1i���N��|8_�<�4l\�Q�15�}���
�-2n!������kn�_6��^l�C�9ܙ-ĩA_V
��s?��бn�g�3wl�y���Ts���XI��>d43��τ��&�E�,B���iѱ1�7�vJr����61W�-��%�ճ��E�XG�L;YE�J~̅��}�Go���ыc6]0[�ɶ
+�/�6N`?]���̘Gfۜ�A��@r�r���
Zݽ�1�kY@2��YԖ��7W�QziB5x+r�������j��8�f��D�2�AR�xw�7�<���Ў�
LϷcs�U�g^���Y���ER�>��ip��6@x�'�h���+]��TM6όO�_2�`o�C�O�>�\���	*�J搷Қv�拭�`s���?� o��3b^ᖻ�&"@�(p����`p-O��p�8��t`��B����ӪPnk����	���q��Q��D�؆��>n.�۪8�`�=�ZQ�S���A~\"�y�ta��������a�6=1j:��͖p;=5I��O7>CY��N�.�7v����ɹ-��)�3��ƱU����~��}T�57P�2�\V�����K~~�;YR��[����d�iMD,̪B���\�����O`�<~O�wQ���Z�b6���"�n���c
�2D%�% ����������{�0ߨm>�|����������u04�<�^Q�+�Ij����jbb�SÞߊJ��=)�4��0�M	ʻd��nc��N2�	e�/�s��4~����R6-U�� �x��  4�)�I'&mAq�q-�8P>��"���ѻ�_�>*?��F v��lRޝ,���L�!�rQB��b�[��_�U���E[s"�y_)��z94@jH���"�m:��]�^;$��RB���y51�_��0G�# ���$`��7W6A�U��� ��X��R���v꽩=&,v�u��u4)�9��}x.n%��Q/��NK���$�H�n ���C���W�B���Nx��T�ꊥ*�����<�rak�a��1D��@�/X����L�����c������z($��L!~'���3�뀓�٭)��ߌ2dΜ�Ǜ�3�p?ݩ���Y[jH:;X�8�e�Q�T�P��vT�s<N���@���/Ј됡+�Լ�=W����p��Xa�!l<x�[Y�#4F�)YC��IބX��W1 �:��u�\��DЬF^~垉!�����=���1�m��:'�CC�v��H�=����pCi�j4��nr���&�Vݽ�9|@����'����A����-T'�Bv���P��]����������e2T���y�'Տ�܏xna#�#���2�G�dT&���OPShk��/P �#̷��������k~��j7�H��h#�I��S/�����FrM��	{=�q-�=`Z4}���N�`�\�0�>�8�jc�*��B�\Ѹc�y�^L<1��I�[�ˎ���t�~Vo���iy��%���"����9��2��\����-L�u� 9J�n{�=�ϳ}���Pmϭ�rVʿ����i�0��5����B� ��A�î�Z�����a��`�rǛx�xF,�<���]�����0��z�wbRx´[JS	�4�ѯ6t�fo����42�VIY�����V��M3	9�Az�P6C	��0��k�[T��%оp��Z�m��3Jsa�DH����jY���^C���)�^�L�"���1�'|ui�� ,|��p(�9�@<��v�	���=U6����菇)}]�F`� ��^S&��۽���J #bVǞ�n��=�õ�y�DY"�Y��=�� 61�!u�1�7;�	\1Tc}���C)�8�C ����+����v��kG�ɳ��܆jv��$Z��A�.G��5ʭ<�E����!�� �a�o��!�Rߞ�L�}L9�/��ݳ�B�5՛:��1|JD��1�O��>@�ݷ�YF�Lp�1[���y�D�T96Y����^T�>'�� p��~�8^X�^F���l�0���"{M���|v4K���A2T���S�]��/g��w�@qrQ�c�n���|����vxӏ�E �3'�O19p��^�a�c�K���;R;���`r�Z�[d	�@{��Y=+���tԉy�H ���ǉ{p"�_C}�����"n6�	�@Lco�X2�c
�T�-@��3PA8T��h�m�y��WA���C	5	�1%�\��.��bs��)Ϙ�?�*P�"=�|N��v����ۛZ�.�����/�H`�����
�|����)h��q���2*"@U�P��x��,�fB��|�=sg>S�0A��Z����
�#J۝��\@��é,E(7�3������7��k�`	*ӟd�k�F\R:cyߌ@��x�I����B�r�k�PUJ,`m��~�jwU2�W���FR8#~�^��.�z>(����܅�0`#���mR.v��E��Xu@�K[��������5������R��I��^3���Io�\�o=�a^\��A)��I�	���}+ ���8�O��3bs8��:�Y���St�s��h�9i;n����7�^��M8�#���ROg��^��k�\+���h���Ϳ������%�' ��Q��sv��W3soxo}­���O
>���q?y����#ˬX0�9J�[��s�.��0>
Y%,�C]��"bp'���|ei�`��9v<v�'
6�؈耥�߀�/@|�B[N@��)Η�$:`�N~�D9n�T��F����;�gA��kX��]�݁� e���N�\2|kϱ�ᘃ
�q~9����핫�.��e	c��?	fJ���z����6��Tj}��x��-��qgCI.��b#��E�f�/7���`����,�j�,FR�2����Fo6s���v��4�v�qg14�$���Dy�Oܺ��z��6�`?�uV;^�0�y�}��"y�'��Hw-{�_k�1�T�"k�bUg�}��CY^�!�l��J�?G��W���YZ�h�6x0�Wp�8����m��W�y���~�d��ͺ�6��^��M� ��)	��j�ȸy��R/,(�ՙF��[g�)?�&� ��iG��U�^�'ı5ӟz��W�P�28�}�U��,(�#3��7-��wʡ��1y2�ާ���{�졔-@��Gy����u�y�c�_@�3���A�o.�7���c͠?�oSv��;j�1bƀ �j�X#5(���cqNŎ<I��$�)ܾ��}ף�����rd'�k@k"a���-�Oh�Zn|u8m��}T2%�|1�AX��c:ݙf+�O=�����p��2���}��4�)��k�J��ظZ�ʨR����->�Yo�X��݁�\-�Re��lךH�(�M�v�
$ .mo��5}+��<��ۥ����tI�`��^b�#	��G����룙�m�_��k�#+����y�b�s_���'�QI;�p aO4ʽN�ܦ�͓b�L�Z+ �^���s,.���3H��+;�M��S6��Z%G�U�b,gH˕W�#2Q����Á�v�� ����Lž1�QQ[�b�[M8�:��&�������a�_�f��HzxIw�^I�͂���rS���Q�ƳڟGa8 �~W���3����*f�NWY�
��_@5�J�븬�,�U���>b�Um}3�;�����Q�i�A��:�߇�^�s�J�:0���i�L��W~�A��q!(��s&�?�n�^<ɶ�����Z�#շ����O�z��q
6�)0�{c��\�+c�νm��^���þs
 �S������K6-/n��1l�<�z��e�0��%��Ygw�\"�F��[e����9.뜮t��(F�O�Dտ�ɜ�!(>lO�A�����l��!&�qf�Z�Nq)���iP=��-��i�!����/'؂�<_?ٖ���M��� ]����$	l
CP����0|��~:u�k�h����e5/EW��>ٳ���α�.����<�s�s{� 8��H^�+`��Jϡ`mn�R~! ��X��ꛔ�������N�>�N�֦�_[*kbW�X�.���������ǲv�P�%#��(�0P C?�!�;�=�_ߤ�~�ku��1An?4ш"I��:'@��ú�s�?o(ѨLmE	9+�%C�RΚI�h��|�DЏ��|�PmykEL��a�����!f���V/��t�qi��WTz��^�v溤�:SLXм�\D��ץ8L&^�l�����ٳ��Ĵ �N�~�n[]L����DІ�J����_��(Fp�"�,���~����L��ּ�����tR��F�hpB�>�Yvn��(t��=]//��n���%f�O �}eu>���]x[LzԖ��� ���n�]a��^HD痘�	����ޙN�j���m%[��
�'Fܶ}1ъ��J���M�Jc|H�_-�Z{�Hg�����x�'Q.�Mu��k�a� �d&�:$Y�&E/$�-�2��ó\��A�i��C�J
���\6~c�k�pF�=i��TD	�dU�8�+��ASb�p�6���Ƒ�ѭ�9⌃k8�4E�2�4jQ�	cq�-n�	M�tB�?��1m�x������F�C{��F�g�k2��S*O,�vbT8px��|�m�T?�c^��W�p��K�vOG����
���ڧ�e	ThSy�e�/	�9���.ۉm|�:r
��|�h�����q���`y*��}��Yp(ṕ}�y���ϔ3t��U[d+(շ�Y�s'W>�i��IX���Eq�L���d*}5�xG}y�����꒗��kD�]vwvu.��>T��AZ�!<�����y���K�&�Y�ͳ �b���CV���T��Ӊ�ؘ��G�h��Y�|�]�43 ���a
����<�R}�����_В�1��wm"	���W��^��t�1g�-KԹR�?b�����y�Y#��Vӫ�C��L�Rϑ�Bz,�,��n6����(�||,i#��/3��f �{��J,�5��N��fE~�1�e��U�R5ic�*����X�k�1��5'�ӥH�	yq\���	���6�ӯ�Ȏ�|�D#���e����S%�&�@�^-)I��E����fzM�gj��J�����:$��R1�|f�Yb1�tH%ݠ�]3�{ر]�Z踽#H[~f%
ߝ8�^J˝{���ۿ*ަ̬3J�<w����%	ӛ��u��xi9�,lE�[�Ĩ�7��5C�ǎ����TU��w�,�lw�R��.:�
90>D�I��~�2��"�4mg/A��ů���dH\�cO�I�t�ު�J#{V#Ș�����->`���,t����UE����ژ��,���B����GZ�:��2>O�mE�6	�>R
(h�e�/�;z)ISB��>�0pʸ��ԕ�)9�o��i��J��"����c�	�UڏؘÙs�B[��z����8��mP嘎<�8j2#([��/.��6�]/�Q���s�O��?a�2���Y6u�[ҫ��!����-+G��hV@�2��~5w^)��V_]�s�QE������Ν�����d&��W���Y��:O����d���a��f>���a\n:DL?e�E��7�hy�`�;�I�έV�e�B���b����@ݛ���cB*T�o(.�ܴ�d�x��5J������h�d�K9/���R�O��W"=ϗ�S�.�<�����H��/��#�-;8-��}`R�MZ��w�����K7�!`ũ�������`4�S�6�+7�^��:x� ���`h��Q_j�ELΝ��	`'������
hzVN�P��s3�W��/�}TyI@..]-�����Q�3W�|�
���� 5���.�Af�����޿���+fk�Y4H ��Ǽ��H�w���M��s_�y�9����$��̚�d�}�}����g���GT0fk����\�`�zc�]{�ߺ�:�p���_�qv�~�z��6w��*�.^�A��Mx��X{�h�-~���Pc�$p�(��⸄?Uj�V؛�ɵ�"�!��E�*��:
�LX��l�U[j��joC=t�J8W�-�9���5f���*e�R�����d;Fg�B��Wׇ����8Twn!%e�����G�`&W2�\P�ٜ�%���qZZkRl/ðu�r��5G�7M�ʜ�PO�g?j�D$9�k�<�^?��C�+d�5�Ξs�w����6�~������f-�;��Ͼ�i.�lR�ztw?#P�q4r}!q����E�>5�m��d0cu���Mxx!©k��ApɐD	��H��������|�ۉ�� 1w(�]zm��{�O1��|��)�KG��v�ɸ��":��d�gE�L�����|�D�f�{۴]/�L���8��엹���*�u�̵��~�U�=��N���1�C�^��MGZRLL���o>7�K}U�ېw������	]����H}ܷI�pK��TR=�Ju�HxH�`�񇱈�V8p1��'%��V�t��#���]j, �̋�dv�ڂ�H�m�=5=a�qج[��Np�R�����_�NC�J��	�&����!S��F��@B�������\��_�£�hN@mVΕ��q����qÔ�R4.���B�Aq>�W|CuO��&K1��V�m��7.vM/������f���L�ӯ�Dr�k6��2�@�������� �6"p�g4ǉ�b�N^�A{�.�br�C�h��&�����s4�'���;��|�]ɔ�ص�"��2K��D���vN<�v-Z�R�YGsLK�%�<2lAS��)|���P�[�0�q�t���S��W*���D�-���s���L�VSZ!&}?���e��F�Y� ֨j7���'�جցJ�4w0��1���N� 8��}��@w�fx�g�� k��>u�*S���B�1�bY��+
qz�l��ۥ�w�'OG�BtӾ��d\Q]/���F�ch��p�r�$q3�!v_=d��
�(g��	k�ģf�!#~"_:�_��L;{g*/��嘿�B����<�}��M+b���N
��S�����]�M ����/19ɕ/P#�{;�-n������M�_K�l�6�g���"iU���j/�
.f�[;� S�#��� j�XJ�CZ	y�*��š����_f�r��]��6���5�9Ɛ9gc�Q�W�JǙ-�=⚹�
9����&u��[�
oL�p�}&����/��0�+w�����ڣc�i�*��Do��V�h�]c˻����;���p���Q ��`Ɉ���~w曥7�ɝ| ~����˿Ct���+7�j@:3G�@�jK���2'��!<>�x�3C��� e+��?��m�.U���J{GX��7�@,����O�v�c��E�]!ȶ�&�7�җjx�abYH|�x}9Q�Ȱܔ5��ʨO}�� N#�I��v����컓T�og!E{*���QP��Z�0D	��&Ɩ#6�e�=� �mQ2S|�Ϣ[ K�Xv��(K,C��Ӱ��DD<�\�g���T�ڦ`�����Ic\mK SFDB ���w��DS� ���hL���#β6��g�)8�erbQ��ύ(���.A�D7��9���q��+�X� W��ߴ�{����A��h��:dj����wq�Ӊ�&֎Luz�R�����L�?��;��O�%��)&�&�Ak20��ц��SrrTHp�Qޒzm��7��v"��D�Ņ���_�yX*��)cal3PĖKA��K�_��u�W�@�Q��[��u�~��l��eh��|L9S|�:���;��5�9]��J�%W�䂸3�S�D�&1"�'�\�+��ϒ�0\�X�#ꢨ5�N�0196�r������u>k!�O8��E(!���0�Sǔr�YA��	J��GB�"z��1��)H����lU�"�@�f�<+&N�Q��P@^���֊����h��0˕�1�|�a�ʧB�G�����F��؝�;_gc�Ӱ�p$�I�C���S�h'���+p�CY����ʃ�p�L���G���µ%��В���mA�9�]{�m:���31̧%Z��G�5���QHv�ѐ�S���<6ˆ�GТ�1 �*51���su����ޒ�S�Y�=Y��[��v%��r���d%��\1*�@���.�W�uO%��Zۗt��\{C�P�9c�w�cݳ�H#EIwH�{���лŭ��/��CS���;���Խ�e�֘�I�����䫃t'F�v(��	W�G{p��=�5�D�����R�c�R�>|�,�!8�h��+�� EA��)Ӿ�����KVs��C2��QHfnJ��׉`��`� �?����:�/����({��@�^ȷ���,�0*ݺ�sz��;��Ug��|�jY�zﱶ�xna��R���f}ے�'+�o�t�yD��@��a�"�ι�7˯#�,��x�ܤ�p H�>~�nUk�f�����@kϹ�A��F
I����	#T�Z�R�����.7�꥓f�h~�3m���"P�p��g�$+*W[-F���H߽�� ՘�&��b��`���v�)8En�S��L��&���h��6!]zc��:�8v��w1�쟸�N�.�{v�s�j�060��M����x*�W�%5����
�_膽�{|.� &ْ�B�\��`�k��qtR����	'����_���4Q��*=����'�F�|b��E���ȍ��'
�*U*H��D$�;6S��$�̎�P�UA�z�L���͐j�5�Ч���h������?.UM��%���i�^mB�7G`�C�
@�,®qne����x� ��y�mbЕ�&�E9 >���c��L��:G87Fm���)�Ng�P�F�Y�)$�b@���`d�� ˂j��y>�/���W۱P�u0s�$2�r�,K'�P|�y\h����Q��t����J��m�9پ�´eq���p/;0S�٪
"��!tM�2�����X��$�[���*D����h\Y�|M�R1�%=�RdȐ��TK!�*y��=�P��J#�\wR����@8`�7�v�P�^��+�]£�H�Í��#���v�x@b�?nmq�������-�b���Aa�˘8�b�V�S6!X���8��M�$�:Uzm/!�.�8x5��>�#SLQ�W3"cJ(k�8N�D�t�;\�F��u�#E����G�*�l�gG��=����cV
��M��Eg�ށ��cq�9W 61��|d��Cv8&,4�C�	��'��������W����?�^\�t�du��g�����R´=H�Af
�����퓱��W<ϠW=2/�S�`��g�j�z)������f74΀����v����R0�u��{�`x�P��E]]���e��@ܵB֨�;�;�\z2�oϿ~�v���(���E����_,��o̟r�IWL��%�%� ����6�e�$�	���a)��S����ԫ�\߾�(SM�/�9Jw5%DPj�@k�u�e�|�"�6���rO�O�K�+^��noM���¶+��sp�*�r����6<\��~��Uh�DXR�sfNC��y�7o�ܩ����9é,C��u���|1'�QL�Br��)Q�A�:��e�������e�p�Xl��f9���h�%�"�̩'�0�8c��-�vہ�҈K_�~��i�['�
�\�C�e��@}h����׏ͷ���=3�������߾���
+�q���e��-1��N��d��i��w]�Î�{𚒻��(ub�[�c���lc���\��^�0�������P������?��cP�4r]@_MzȻL�q.�B�G\��3~��nğ��T�( {ϷM��*���pDwI��X�-뜳��tK��pS-��������m�����g?��zm�z-�<EqD� 6�M@?o7cT\�٫ 6�k%��X3�i�i��f��QN����S�m�e:'e��[�D�M"_4���w�!�U�Ma5�3k�b�-~�Jv-5�2N�R�[Q@k�m3��!U�fF��{��"-��#iHm��n�|�fx}�{��'��-%�Z� ;�%G�W� J��wKW�X"��2j�BX�2�/y����Y�N\nqЈ�7^D݅�cE�qY����{P_XۭKnnjm�M,p�/�͐��?=�k_u)Ń��~p��?��lQ���)��6w��H�d��,���F���|�����i����C�S������`A}7(~��8[�疒�����ۤ���D��<���1zq���j9�HO���2<\{M���s���PY�Eڔ���*�U���Va��Bxe�9�p�.�����P@��15��;�`/��_��'���!�3����>�/%D��/P�x�1ji��2>���Rs%[#�'G.�pPx���^�K�󑔚�v8��>�es;�]�Z�2�1�9��5Z��J1�k.�s|��
��h[���ե�L�LA��X�=���H�[�:�0�ǘH�&y���R?@�c%	s)|r�֫�.��PF��{�^4�P3�pSU��a䬣������W���в�d��fV�Io�J�h,��2�ͲYmVMo��{�)N%�@��Y�����o�Y-j�Rg���X�5�뱁���8n��>��\��˸�A�Eѿ8���D|+M&�4W��P����S��q�s<�����䘐�+]jhgg�t�<L�)�u��[ڇ
"�M������"*P�m����'yzL�sv%��ľ����:��^wZu��
��$V3\@�Ʈ�1�В/����G��Z ��y�ӷ8�t<��J�Hr>�w!���Uj�<X��TK)ѫ��H]���m���W{�W5����ۈ��N2ы:�>~�j"UL~��`Eʅ~�����_��,&U]�>�����u-p�N�k#�lu���E��a7���_) D) ��@6��=G�IU/��<��1��X�:4B�2@Vgw�N����yC�!�0)�Eᑬ"��(�Mx��0��q`X��$Έh5�3�z+  ��g.h����n��or�4�P�XH��Z�4���cJi���ZA�!K�v�@�x��˼�e�sX)���Aeȉ���}��K:"�V��_�aX��>
l>e�	�Y�M�M8(�54Ig�訡Fh�6���ڤ|؍o�A�-C�. a���O<�S%�y�zɯ��C���	@w���/Z�s�3@�5���"~�Xp��Ҏw1�g�F�Ud� D����ni%�p"�G����ؓ���й"�J�����1�_;K�b�U�C�<���'j�4��<K'��3�)���D���Zח,�2���J_xDU&d�3J��(������I�z�+,�I9j��`Y�������v�&�M�����SNT0�h�*2(Y¶�g����?n���6�*��k�;\̚�C$���o���S~�hUf٥z�����}��h�Z�<U�2��0�;/Ɂ�[��&��l���e/ޞ��_�"��5�?�Hr
�<��~�*u���>?���	oyT��fώ�l%��<�[��U	����O+*\�!���"p�6N��A���XtK�F�|J���W�w�񒪵�� ���>�?�A��v)!�l��(9��3�p���ġ��2�U/��������m�?x��%���X��4�h���	Ov}A�/~=M*)e�2���
�S�Y��7m�z��c��Jr'�>�_�d�����������1�ل�2���Zs�C�٠z�HXi?'��8`t	cI!	�v�KZ�1�����VW�y�+=ANR�{��Sv��a�D�� ����+�ǧe����x؈Zb+P������}�`��x����J��w����#́|�)�C�_����|tr)����MX�̀��S�*d���磻�:�ꖠ�*X[��Gn4Üp[��-���7�撝5Y����~������
@�h�࡯�d�x1�V$R��1s��1 �;1�5ͥC�4�}�oƠ�eS���F@8x�������0K����c9��3���\�p�2�)SmO��xc�Xh׌����N�/�	{�Kj�(��+�a:R��[��7~�򥪓N��^~#-^{��`(
T��?U9�0ur�k�v��B�cQ$��SF0c~6ع���' q�z9�Ɵ�.�����l^	�H�	gΠs��»�Kl4v�z��!����椛z̫@V8�z�H�˦��md��� ,ˆ%r��g�n�^���oz��cF���m�D�`9�giX�B��3\1Fw��ߑ���܆�t,��i�i�.>C��c	�1�<�%2ol�Gc,-�$�V8���E7M{�?�n.��N:�Jʎ(�Xw�����d{�uZr��DHOޢ��b�@@����z�,�A�؀P�x��v���z��U����7ε8e�kڎC��h��el�GJ���+:��t5�`50��'<��� �����}�n�[����lo��>�a=��h�K�"�W8{u�~��בs���1�	��"f�I�Rdj�o.���T'�����N�ķi��F:S�"i3�%Gt�^�yzٲ�M{&p��kug��c���9?��3���3u��n'~Ru$VzIA�ߘ!��ߥ��ߍŇ >b�H����|T䞜i�
/�'n:OHî�H��'�$�zx_���\Yk��d/����\�gO)��%�n�9�!v���%��h����vF���e~�㬞�ܟN@��]���C�4K)��#,֛��i�;���Kd��Vp�4��	�����A�f��c��fw��>��Ւ����+۲dz��W�Uߤ�z�P����J�pi�b[柲�9�S���q��� �9�����~^~�7~Aa�P"Zb cw�,ԍE`����ws�9��� ��� �|�-;AI~��XQl/��R�؁�D����6&�;_!:���v֢ݎt�8x�qA�����1
!-(��}�W1��=4AYP&��qI.���@��K�D9c��6T�c��P��~��w����
tM��ir�U_�Si������uܵ��*�E�փ�wq5
�'?^���=M[l8�)��KSo�[BN�L��S�#i��r�ʠ���6�*��`eJ1�:�z�W�Q�ŏ[1��OM��n�^a��n��!!��d`�j�C)���7��~�C�&w������խ�A�]�#^N��v�khO��` Rk}5�֦F���i��y��s���rb9Z:Mܸ��U��#���7�xtƶ9��%��^�����I�4��@ﮍo��ِ��j�	���%�P�V���gk1���Z��e�o��޹��nʋ�x��Ǚ@/�Jk�f���=����m+˥�E
I�W�'�x��()٫JW�� M�$� h���>��"��98�M9a\���
E\���,r۷~��h*5����G)��<L���q�fZ�z��������~��&,r���.���'J��ÝHU�"#jv,�:�WY1i�>�GF��.���SX�5Aׯ���eF����_���t��V��izܹ��#s�af;���m�hێ~=9��,�����~��v,?���TR���c[r��P��]�̄�|]�?SxB��,���u��6�ߢ!�8��Phr)n>��"�pg-�f}��x�� ��ݥ�Y`�D�h!�Loo��0J^�yϢ�.l��m���G[}s<A�r��q#6q��"~?��Y�����H��閮I�䮐(��X�ӯ4��{I��&��y�߾�t8"�s�M�ƢY�b(���r��r�qa�zVR���G�� ����Ҵ0�T�G#��ǯjE6��h^gm�=������J�z��Fn�6\i�j6�S�����EJ��K�R@ɯ̙�W��}/v��0�W4l��)ŏ�h�wQ}�=��`��K��h$Ap	^�T�衫쒼�~&z~�;��P)���Hӳ�0��Y�r���@z	�h������\ψ�_�Oκ�t!�9�����-0���x���D�xj!��Z^���1��()9�}��mP�.t���Ѻ0�.y���O9��R�F����\
���0ʉ�ʭ�=���V}*;��~a�Jߋ\,��8�J�ᅫ�I��� ntn An[/t.�����#8dp~⒚A����AW�\d�6� 𰝽cxz>�#�׵�8��	�`���Qʋ���)�)��T�W��GK��L�V��9��t�Y�_�b��Ə|��%S�?�^�+�m�0������Q8����P`3�h�%��1�h��cF�v�!Ftz�3-�%>Ҩ&�j=$��U�<W�;]1Q���X��L�I������o�'w�W�x�50Ƿ�_�&��?�����7�t�w��"g����uHި�C�մ���U��^Iq����%f�:8^�Z��2{�x���?���Q�J�]�a?0�����ߖ�M��hU��� �V��DW�{���rWmA���P������PMx�)f1z]�pV��q��s�F4 ڣR��!�۪�C�����0�!���"�����;�%�L�_�]o����e���Q���ǰ��4��.EE/��`�0�3�d�����q��`P�z���x���1��K�]xr:s�IaA��A����m��s%��P��g���ހT-�ܚ�&u�ywL��5�!��=����0)���r"�����.H��M�z·�D�E�3D��J�7�����#��p�����"i��mN���@i���mD�t.���~���6���@�0��d�T�<��B~��F�x��i�#�����`O	�Ixip�تG�b���ꦣ��C��;i {���ۗ�?��%�&Y��(o�P�-��g������O�ŀ���'Ec5/k���.�Yy�W�0b<\������`����n�l#n��E��d$�j��1�f!-���S�Ms?)��φ��%��8�v�h7~o��x9���m�m���s���uSHh�>��z�2y�O�㖜������tt��[y��Y���v�HcJX[�eޥ�_���as��L9��wG4hd�'�f� r譵����rP����S8�޾܇��9%V�Y&�!���x���'-Dg'�J�Y_��A��HC��w�9,��ʉ�m]�3â8������F+�j�����%T����_'�-^+�އ��^$�n)G�-��#��� :Ԛ��SX��;�ŋΎ�:���bƙ�[j�����%'0Yr�g�� {�R1��y��vn�پHS�o��T��r`k��Q�5>֛砝�����>K��*�������k5�dNѩ�c�L�1�E|����u �&��\TSy�دh~�l ���IZ�[V ��oZg���ܣ�/����v��Z�^�I�	�ſ�E�(�A�xf�
�"B&KP��)oi���؁���If��g�5F�1ˁ���fّ�1�;�Ah��� k��#.��t����t����Ӄ�9{$����{8t��S��D`"�>�����(��$[�!Z+
�5��D�s�૟�RAf�F>���}	�!������_�x}ؑӴ��ɢ?l߮��EO%R�������$���!�d�
�dt��U_�>��_[á'�U��P���wK`n�� ^�.�X�)B���zrw{���F�C�h���̟�d��&��t��W�~���x8�;D��j9��:�8Ւ�Μ��t��5��+�!�0�����>�,�ͺ��c���F��f��@J߾����T�W�<�����zTbnzDp3q�P�
/�ܶ��9��ջ��ʜS�kT�T(۷�#����v*���/��7�(�M1���,�U2m��پ�:9�^/Ai������Cw��x�7�7�6��$}�Z�VX �|U9J޹)P�&����wwL�~�_�8�F4�R6~+H��mm�^� �Gs�ة��+�B�iI�R*�H�K�, ��t�n+A��t��d�Ţj��gZ���j�����0Gmx[��KG�U�*��Y ��ޮ~-|X��q����%���	���9����n�^��:>�5�
f�QS1;���'3W�&�I3�~ 9�&��&���$���fL��y�� <��x�<�]������@���[~�Gn&��b8�-1�ф}Ubn2�Nߪ���y-F�I��c��z\]��3�+~K��o	���� ���bO�r������1Z����Na4(4odu-j��}8K�f�Z�n,m��"�#I������ߋnfE�sh%jAE�����2�?�(�����@�2V^��,�L��R~k�.ڧn�YR�|vz����0�'�ǆ`5�li�$_�l~ć��`:\/�ble��ǯ�
 ���$�{��`0�����E�Ĩ��	��s��q\61�(���s���d|�O�ܫ��#��}J���	2���[���<��s\��Ѹ)���hqr	=;��ܥt��ѥ�r���2�-��µ�d�0t@�֔m[��V�ן�Z�����?�<���I�����-�4����ɄIZ�`���q��t�}@Q�Ī�� L�+����#�����qd�&�<l;v�I�m>�T~ʲ����9����i܏ E_��"�^;(���W���6K���ܲ�(�'np�y�(�OD��2_���ՇmeJ*ӧ��Mj;H�v�>W!��u芮��Q�`�U8ׅ�az���oK�!�x�6�N,z�^}��6�nqd`�p��R1V�tO������X|㺨��^>�$�2ΩT>y��!�%((�D��A��>�8CU�f��h�e�Z07���I����@�eֺ����>5�˸[�UH˥�S���W�i��-�}�o��2g�&|�1^/�)C���#�*&_,+;�թaAv�td쐂}ς8E�U���<�^��4s����p��L���6߹s/���ce02<{���2�;���H��Zpf	�v����XA���1Q��{��h>����J3Ԛ���q�	���L;��ЎF!����G���p�"-�������(dxE�wz|H�8�pa�x�L�4O�/��o���Y�'�2Bc��	 A!���H%�ք��~B��Ty��.,٨!��ɹ�Q(�X�`��?����e����>d+�c�������0�#(��;��&
a"*����,��/�HqTTSڏ᱖7�
]P�S�S��^��2%|�> F�ՙi�3���?��:&y��f˷�ʦ��ɜ&J#��
�'����:P&�	h����RO5�ӎ���Sd��x��S�}q��v������xs#�[��ךd{`�cm�{O	+�<;/��7JDF7_Ƀ
�R�7�S</d1�75\�H �Ƀ^�ms<S���$>Q:��.~������I$B���D�}JZ����H��xU��*	�'A:�ךf��W\[��ZU��R2��L��f�!��OPE�?k�'�3�����Cqk�fP�ۡѱ [�ڧ����4?d��m�6�مh��ܹ���������3��ͻ尴��Y3�n���2�iJע���~�9@��B��P5�2��L3(.}3��$든WO�b�1�K��|8�q|��)��j�k�6��vuכ�������\;B Wh�E7!��@M"�:��U��4/j`1%�ކ�N���S��0�ȧ����m�����K(��վ��^ �Ap��^������9��n^�!�%C�� Zz�h Bl#��ʥ{d'V���d��7��Qu����T��:٭`��\y6���L�-C�nQ�	"�3����8�m涰����(+��!�d/���+z�<��;���Z���`���	,��Wr��H=l�,D��CX5�ˇ�x�Q`�7S
��%����Si��\>�n�����N�h����8�;�L��3�
�_��RU�/|�.�Gn0���szU?_0pY�t.���0�޴B��ImC����|�H%SCED	Y��9]��v��<����J�`H�`��n�����������͚�D_j��{v����)����^~�wJ��ũD#����{�52��އ�_18����4?���@�=u[�->Ё�U%���T��\��{�����r8��G����0$��St�G_n���[�m������.�C���]�����;}�vކP?����-\].��mE��4	0�ˣ�"������5�+� y*��(-�
�Fm��܃�.��%ma�v������g�ˎF���=��w/z�,�} ��i=��6#� �
�K����7+������D���B�Og�H`ۋ�Ġ��ɼ?��h��J�T</;V$]Y���u�]��r0=�x�y��p�#������{"
�2N�d��e�b>�9n+ݲ/���ԿЯ%H�c��ub{G_<��;�)��(n_~xuPe[�I>�s�k��bmʾ~�tD��M!�~K�Ez�/��m5 "#&M!��懠��������'�C��d^�	��XR9��zE@]eO	�Ժ���L���H��|ڻ�H�1ZN�U�|����z/��4�Q���\�~)l��9�����N6�Y�?]�΂�Z�������f�����W8����Ȏ�QEet:sq�'�J!9:<���$��r�7ũ��:�<�ŏ\�[�
��woX���S�#m�0<g�E��,#�9U���(�WM��5'�����"S�+	Л�rA I����i���a02�f� �=�+����7�ż��p��BY��o7�+�L�M �\�Cf�&C ����]��5B�=�֘�� 8�mᏆ_G%d5Ww�P.����'AU�]	vO��L�4390
.��L/H���"Tm��;��=D0	-9����7��F�A{�l�W����hB�j���@���p���*}C�wG���}L�9�f�\�ɞN�����b��0���q���Lg��l��rϡ�0���}.U�����/�	�B�T�^w�(�kg����'E��O>� Ve2�ߚjr|���k����[C���$ؚQ��&Ճ���	KA*Vq��4��H��i�l|�GĿ��O�������q�@�o��C�}j'e.�/_&-⭃�h�&���^|�ћ 8x�ai�e�NL�Vx���@�-�����������3����O'���H:�l^z�$�B}���2��L6��P�*�F-�v 0*OƤo�A�e���D�&s��;HLt��G�m)Ci�NhI٩��B�[�+3Q�<�n
��Y�-�����[�_�A��=y������o]k5�p�ώ���s�L����
'.9�GȤ��.�h��!�X�0����U�U��D�DR����Cᭃ�$���B�RM�Uî����2e�Ł"�t�Sߡ$a1����!��W~Tј�NO���#���J���׊"fǞ��d>w�1��T��jaU�Tj�P���O�s��Z6��
5�18o���]��1��>�F�@�y#+x��-�DN	�q�7(
#�[����uuN���ƈ��Q�_jfh3��g�*���=;�6K�,�!2=K�4� b��*C�h���e�Ja�X�]�4���X,E;I$�.x�T���!�?�O夣�?��ٸ��	�oC�����U���3��6;�#���J�$��r^�"V�5�wɎl]�\��R.D�W���p�<юX��8+G_v���M6�Xm_�L��3�����FRo.-y2��sa�"V�ݚ7�޹�NlX3=m"ŚI���ز�(��)
wikh���jT�{��? 'Y.=�������ǋXo��]�3�S�Sؒ�T�,G�B���1�6w½+�|6�.F[���CU J�}x�{
`�}��,\B@!9�D�<�%��}�6|�GlϮ��a���2/�T]��}�>l�C*I����C��P�b��)Y�\�^�Ԣ �%��I��������~�S]$��&f���y���k�B9����N����'���ugH)t��0�t��Ô����Pi��fί�P6
��V��I��5Oj[t9��ο�Ū`l��	��7��T=E�.A�{�h�;� �z��N�����36|_��tA���2
���|<	,���.���taQ�G9R1�k�񓡯s"} h�=���l�Z���*2v���D���?��ψ�����?��_�+��H֬;/!E��@��AzFF!�H�go�Y}-�%�u�ЊuZc�4��"�
Wa8�vk��0��{�Q�lOg�X��e��"h� �
��>�A�)��@��-=�s����Ɍw)WEF���VE*�f:M)ضr�j�����4����aN��I�lQ����f2E�Gj���Y���'��qY1�#P�|S鉓�1]Ko�짅��J%Ƅ�4a�a�\�Pv��G��#�+�_K�h��d*�r�-�Y�!W����5��6-��ku�P�&����Ѡ�0� Fzщ�
8 �1q��([���K2S�\��G9��A�Q�-�P��VU���3r?��~§?�'	!�23��F�~�pG�����n��� ����ME
��?�L�zd�Y��ȌB�G�,#k������1Ĕ�u��Q6*�����|��3�>-��n3�`t��-S,hk�Ur7^�X!	���qR���T�y�3y�y�΅��P;<B�|H�Ca�?��Ax�y��8g�D%EY�W'��N;S B�o+
nJ5;�s�r�=�7j��w��H�b$ݸc\f���ɰ�8}�!�{y�j,Ǆ��ե���ݒ|��<�ؾ[!20��� d����o��aT����g�ڬE+�B;���i�:}$wo�-�\W>�Y_��C�|������&/ ��,��9~�F@��OXKW�ˉ6#�$t�����V��|�@9*A:[�����Oޛ��	�� ��[��NTI{p�A�:��g>P pu���,��h�ܳ*s��
�����Es�u��?�`��m-����L$4��T�5��r5u�;[�4�Q�G	TT�����eI��g ��%D�
�/\�ꙵ��'���6��|� �"m9�q��w��@�@F ;w�}7jڂ�$��e�섞��?I~f}�'�=��tIt�ާ�s#�ݟ���^8� ��[v�l[�����O����:�*�c�d�Q�s��C��:������@տ��@q�h" �;03�K��������?Ѳ�/�� }V��]s��j�n��,x���+]������7�f��F3&ң��`�k�I�����$����r��� �Q��Nvh��i��緺�.�x�h��=Դ��+Y�6~�]b%�^��;�����1�"�qx-���5_�$�T0��k�D!{;s�X[MG�7�8�D���VZ��T��j��z�|_C~SMOezl]���5����x�2��,+�̰Al��&�=� E����Ӟ([c�s�:�H \0��o��ص6��E�,0�-�9���"�JX6AO
ʳ{����I�icqg�1,wۡ�Եd��&���A�d��洧�[���I,H�S=������l���.�J���������O�H��"��t��Ll+� �wW��
���iD��ө��*��,�;��~���������
�3Wr[�q��;��̥K�E�������⯲Y4��>4�̨�n��n��贓gS�f���#uɢ� a�R_�
�QA#J���8�a��ʹ\�O��M!��P��,D��(w�gn�jn���'	�F��U���/��	�w�,.t*����Օ�,.���2�����g��#���dNށO�S�0fl
D	h��'n�����B`ܓFf�ʙ��&#cN�B�	�۠-�(��gM�� =Nx���~����L��;��v�[MB��y�|X0�BL<땒�
9�&���T*α��6^)H�V�PH7�.�i�� �&x�3���,=F��4�ө�Y�ȝ>Bzop:��y�ӱ@�J;��4���j[�_p�����B;ϒ�	�]a�׻l
@��;�o$�Fj��������� ~O�������@��f�mu78/j<���T�TQ��Y�Hշ���yP�7T`��I)�����c˂���qď����&�}��ȥ��uM5A�%�ȏ�7����Jfm +��Z`��ǋj�^#:�)�#�Ub����Ԃ.�:6W��B���`�
�Y{�/�aA�A�x�{є��^e�[틨���,�]��~��^��j2Nȇx�I�䟋��:G:�>���p)�k�)�?Z�Մ<�۠�����t�T�t���"O�ߩ��/�:�P/�ѣ��YY�S�6(f"��G
�m�֩�{v�SD�FW)G����2�jY})���n�k�m����՝tE����b5�ę��ti���{�i���ը;ky!�s1y���%��K���ٽC�)�Mv�{��*�b���i��U�{.̞K��ͺ�`��ʳ��087d� SS��k��50�d7��q'������@)z�����n���a�!�~����<�N��[�=��[y��Z=�J�1+3Q{{9���q����U�5C�!�\q0�\PM��I�M!L(l뉃"�A�v .~8ZC���n���J�k47}��&�h��KJgtsW(c�=�A�	bEoI	��M�t't��:�rcmK-��Z]�#�6���h��N°�!>�RO<�e�Ft�w 9�� ���U�������N�R'(p�d�Õ��p[~�Y��y;k4=��.;^�0��=���W���L�#¢���t?W|x뤅�H�b��Lꋼ �!�!i?�W��$)�9�;�9�s�T�g��#���4�T�  �V���'��>Y��v����V���N^�t�+��[���Z�j=98�aT��VOL3z��r>ʏ�Q�E�rv9P��y���!ɧ)}���z�fB������mp5N��s�(cB��r�I�V�:E�혗�ɐ��NStn��^�u-��2�b<���Đ��Ľaj��}2˛,u�F�Fr,��h�	k��T�26��\.�FtmnR<)X�X��t 8�U�?7�v�+6��N~�7�O �M�tH�%:^��<�����MG�{*�{�U1�;�C
����c����{>���Ȇ q����G«�Р�ӚyM膡W��F-d�
$ܒ#5�/�x���A�nA�x��M<��)HչFw�m�9nP�h�K��h�������$�_>Z�F�λ���F��С���J��Nd�':�yK^o�2���r�M�C���pdf����L���(���ۮ�=ŧF�M&�Lڤ��?u�T�&��z�I�	�0���`��40�?Ύ��@="#�he�Vc���?4#�]CH��H��w{M��
\&>���� �@sP�g:�����f�!v���L;BK�3��q���@�)G�$���k_��_�����}A��q+["=3��.(4����]bU*t/ހ�X��|*�*m��y��ڃV;�:iU��`���������Q�4�Lp�}���s�>Nq�/�Xy^��cĸ�)�����1?��À��_�Zo;>�3o�^��^����ȳH�F��:�]¿u��T�Hu`*��MC�p�+7E�^��۬�-�x�XV�T��s���6G�m��#W��▪��\��;�Ӡ����4,>[lk�������=�G<l&��]�IG����	�׶�>�(��#�\�:�8~q�<�ywm�=1��ӥ����ӌ���7t�I���=�Ԡ��O�B�/Q-��AQ|!B����x���W�N��*�y @$"#������81���=(l�F�i��p� �yLt�C��|� �*��.D�������.w��{��4������i';؂I!��R-�g�6&��ï����6�@���w�um�+�L��~--�v�f��U-F�v���R<�N κ
�>Fs[B��Pf�vP�#宂C� �3c�WF��J�=aR��\��l�;�u�k;����A?#���$ԧ0ِ\F����8])7���%��(���ݹ��|�w�m4��0$&�W���*!;���
�Q�Dc2da3�*��MP�Z�oD�6ķ��X
�`��\���o2�EL��C��#̓(�'(m���^�U�/z��{^��A"&���SЅ/A�-�2~������0XJ>֥밣���!�Ep(ub����*E��5���T;�M�������"���h�z�%�}lR�7�u'c�@�d�=�� (ir���4�EۿB{7��q�x-�N���.�>����陬Ɉr"�6��(A�&�S�\�v�4�I[�����yv}��P��W�d1��_��"��E�9�<D)=���=BX�Җ��%v������Й e��.���"ԃ�B����󳮥Yzp_�O؄�q�2՞������i#���hyL*ݛmuל�LT��u����A�Y[��T"�J�)��L�FQKr���b��D���y�+ʘ�us;q]z�.���[�9�Fm�K'Jv/7�<Q����?�s6$�0�R
p(�v�s\�C`8�ߛ���[Z�@RT��g�Ǣ$	Vj�$�饪��Q��x o���/8]���-o��;g_ �f��7̝�W:j�Lm�$](���`Ӊ��4t=�T�P������r�a�:��w�����݃2�H���B�#��̌'n��4mu�gkN�G�����d�#Ι� �������M�A��>	M��:ہ�;���}����Μ���`l+��?��'���/���ձ��u���0�5at������6�;|�OB�q���tm�2D�A*'�/���f�e��v����T晛o���*v�i�m����ⳛ�n+U�-K�����t�7}c��Gs��M��봕��u� ���L�W�YY��O�:��Y�����Jr0�Vh��DގG�ĭH���8o�v
���t�̀D���N'��*f��F�5��[����(4j� �����l�^og{%��<�H(�2��9��(ه�����j��S�LZ���M81��� �Ӱ��o�I��?�1�yX�p���I���6`kZ��L*�*f-��o�³�I�	ip&3�?<S��Gy�h�16��_^��[��G8�T$�0�o��46���ޯvlE�J\�<+����O�&��K]A���s�܋��~=Ǉ~�ET����!�UprB\�n4�a��q=vK�#�,62"i{{<C�����5 �2q��K�ݻ(�
(����?E-�9(H�@���:�U���_Lg��f�h}nAGu���ޥ���������	k��3A��]�Ld�vt�t���q���z��%G���쁝k����~�7β�z��y�ເ]��� �ׅV���ʅ(��B����ְ��yRK����6��1,"%ǳ;r0B��ӆo��wS���!�7y�˭�ڵ�O���e��Z�ŉ��%��H.5��|��+�� �|=��-$i�Ԛ�@��Np�ӑ�};���I�3(�>�G�ܻ)�`�m·#i>g�7����מ_UT"�	,��|�`�������-�Ȍ"�ӓAF��Ѷ"��P����9�ر��f��o��,\�؆PN��:}<���O�z�|���Q�z��ϐ(r>��c��Ͷ�������3ζ^8wӞ�nN�"H�*����%�Ѥ�Ŗ���ෙ�}��I��-�k����}��']��6�ع&���dO�,&��=�Z,��H4|��� H��i�l�SE�
6��'�V�*Ǝ^��ctZ����W�}��+{�&�|X����y�yM�Q�eu��}<�B�\h�ԍ.ç^������/	�O�sE��bZ�t�-ǩ�U��9E"�;�#���%h���h]��@�T�STLAש�� �S�++�4��^�h��P��f/쮵��+#@�����*X�:#,�4'^2p�L�yQc�"�sڵf�o�o~N��|���-ȭ1Ih�i�z� ��%��-H܌ę�ـ6̲�c�2^�=�ޣ2�j=��D�hg���y���j5O�i/�0͉�t]B�(`3r��{|X�h��	�ǬQ�l�o�R���O��X�\�%�+]�[��8��R5�d��
<6v^�9�|B��k�B�ǎ�q;�9���̷��4$��>^x���1�'�&|	�'����:m	�溶O��0�������k ���e�G�T�^�U�+ܟ��ά�~6h% ���9�Y�?=?��v/h��rxh6��Ɗ2/b�c����]ײ[x8���mZ��s�eP�?�V�����f�q����3bSv���0��Xl���#�2.,=��i~��fA��wԤe�����0���*�4�-�]}���[��9��{�[�F]�����H�t�d &�*@!��=V��Ofeʨ=�X&Qaݱ7�����̨rG�TS:� ���kc����Ե[	�h�G�<�W��������G�"�� f�kى{�J���%_�E7�lo�9��`H4�:�vʄeǩ)��؜"�Wv�D�[q�O��iA{��Ȍ�p<��Z�	ac���)�e"kB���YM����Ƕn6�>�|M