��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�0b�:.}$h�&�+���߶��hEn|-V�d�WC�j�G��9�^9�-G`-�̓@y�T�����d6g2�&�͠b�^�R���MI��s�?Ct�l�����%<^}���;H�z����H�>A�:��.�d����M���P`�����_|F��30��@v=��Q��S'(!`���Z�D/>H���1�s	܁jb�'�)zF���Ƥ��#5-`Bu&��LUT���m�0�M*����uyO��=�_DJUS!(�79���U΂)��X�;�ܠn�.0+BTV��i�(���K�!bGzx�0�,)�']Kxq�=��%C����_e�DP����B=�lW(mQs�r���+Z!���9�2���Бս_P�����EO���䞿��7yt�*0֚���
��z4�RC�AQ�>`���ԗҫ��y6�������HO1��ђp�Y�tGkᒃ�z����W
�p�lAl=s��W^�@���m@m�Z~�YE���-Ƴ��k��Ƥ��D	�B�k�q�'!x�G���+�4\���1/٪#s���<D4��A#6�c���W���0*����etN&�O�l�Ha_��9�$����q�^"�xbyH8��2���9Mg��!x�M-���a���'�bH1t��)[��������xQ�"}��l���F��	WZAc1L �U�lף˥Yth�#�,ыT�Pũ5���*�Ԑ99^�
�Bc+�2�g[���b;�c�_^�Y�y�i�m��J��/"���{ԅ�qI.C�^��*f�Zk1�ds��C�6p��rFI��TXY#�/K�!�f�J+Z?� �@�-�akԯI�� ��̬W2�F�mW�xZ�2"BO�7�75$�����?�ښ��j�[����P�D��� y�?X[]��/�('�v�2Ò���Wg������-�i?� L-�����c���O;Ps��?�:;�ǥH�s��+������g��^���j������n��5[�P�`	�����!wUM�M|�����(���H�N�&-�An�4d�|����}���FW�B�;�s��l���{;Δg���`k�Ϫ��6��dW���"T�0���P]чpG��|����<������"�W21.���q���y6k9W®X��`z��=gY|-�?Mg�³M���ؑ2��n⽃ʫ�x������JNs��터�E	=�`_�( ��;��G�m�)}�6v;��=��I�x�s�jn3���w�2������!�+�K(v�Q�Ⱦrx<{���깏pc^��ەsk%�*���ϙ#5��Qa_�u5�A�r�Ia����j�E$O$&��b��K�ȗ�;+�y&@̟.��a���Hߩ�0����P>i �^3��PaX;8	#�&^������N*j#��,�e�(A|<rV�,���N*|��%q�6�������ڟu�&t���Rzz��Q|t��[nk��� ݭ� ;]8x���l�KQ0S����$f�'?  =�چ���qs(ybZYPe\�4'�;�`��""�0U����nOb�Dv������ Zm�'|�1:GRR���t���Yo�	��ߏf�;�(��T���XD�P�;�\�����p��Г7z�:XG�`�9�dͯ ���1G�����KI�(^��D�B*4��	��+:Ŵ�#�S8Qv����Kǻ�<�]����;<���W���)�CVC��X���� �8�����k���Z�w��y�H|f�8�����!`��QuW����$>�&�%��Gp���Ô�4�����]��  �8��j�_�;a!1�R�����
�9 7h�4��s����7~w���e�o��N�1i�+�k&�fjIHen^Ŝ���$<x����\Ó�djiٸ�^�ث�t��	�����D�As��o�!�����)A�m5�P������u�5����rx��H0K��]�
|�(}�$4o 
��Y��Q�w�����8�H�d���0$.������y M�Cy|RN�ʞ2F��w�i!�����zr����^ 2W��-���6�")����	��g��5��Y8���ۏ7��Ѭ���׹��kP�<I0e�7ZfN#��}E��~.U�b�_ǖ����� ��N�V��?��7n�p%�������f�嗢������~�"��Y�yH�<��o����+�	[��6|(?�C�K~�+�}N]�}	��₸47Q��K��t�?,b�A8��kd� �,Eܴ��~(ͳ�_��������}��sz�X�Ŏ*i����KipaO�>@��I���z;�-�%��G�>rPMq=+!�v�*�7
�H��D�"��ѡ�O�\ ���R~E:�|2�D���&� �^H�xH��B~�}g}�O��BVWC�_)���"<s�b�an|rF����wol��Fz���H�'�)���, _D�U�4�\�Dp��Fu9�H���s�\��%!	�i3�����i;��I H�_�K����xtC�������$��`L��y��_\=��JT_Z� g�ƃ��b9����%��?� �����z��l˃��;-��\����q�������� 6I�� �����ƚ��� ^i+l�r�Om4�}�OE�=��ޓ�o_qjv&!;��ӳA|��e�0{�a�{X��Y��X�aꏱl=�;�߶t��M������ݾ}��5���?�����؈�[�E��,~a*��AN@rQ��O!G���l��l1ϏSK�����J���D���ݼ�V�L?����wIWQ�K&� Z�Q���?,���|Fw�on���<Qsq�\�ێ"�}��{�w��/&�
1�k+��|��2��f�,3�����)�c˨=͗4�X+�����*�X+���p6�H��`H���x�7s+o%�:�(���4�
���y�S#`�QZ����֐6i��;F/z��p�o���;�}S�,�b����L>+\uX�\HN�2@K�c`6u��bJ�n,~�;d~@q��IB:xf��;~:u6�(��>w�gr�E_����`J���q�`�|�9D=H�J������1� ���s�����u�7�<C�=�Қ��2F���2�������i���|��:'��J������gd���g?ѓ*�űC��9�Y
��bIڦG����F�H���=!��Aв�Ұ�V�2�}�􂞧,�z��6+�u|�0�S{;�	�E�?�6�OU s/��{`��/-��S�?����qJ.�.���&�ZVi-EʜA��Ц3��Q1*����Z`%����r̂�(笴	��.ql�3��]%k �rO^[R�;"l޸�$�Xa�\v"�h�(��|�.�a�Iza�Z��ʉe���C�����'T��RZ<�ݬT�J���� �f�y�uJ"��d ��&��`���<í&#�{���x�Bn�"�°I���U�����!��q�?-*�IS��ge����]N�`x�.�v/"|q0���c�:6|� �2�c��">��4a���ݿu�Dٟ!�

��&KOK�2���U*�f({��
���( cjw�f�&���5��0iB��A���(�@���S�v�)�}�䢙�vNU
+��Z�������Kn}%J�W�;���('l:iM��\dfI&2=q���+���s$W<���;E�
��O�+>E�F/(e��u�N*�$���5���\D��xTH��v�Tyf� %�6�BA��ۀ����5��g�O�S�Nf�##7V�+l��o��;w��;����P�5�ڒ��:��y�+�|?�p'�)Z�r���V�dh_���6~�Uυ~.���<�ȟ���V��ΐ�.$y�yo��*�����!���VQi��m�&����c"~E��)�И���U��'"�V[H�-�����@��m��ųd+�ٕ�3��p������v���n��ŤH��T
���h���۫=����>k�g�)e�XT����t�k�:3���k��e����]�:����I��t*/R��:�7�D_��8���-|�<�16n9�[�@��ХT�5���!��Ė����O퇊�7�Їۃ�!jr��&���>�f!�Hr�:M��[?��H5L^h�� �܎Xz)H���'���#�;1�7:v,|D��$�����BI���C�nE��e� �l����j_) F��g��z�spF�l"��2��#W�$�JI����tV�ii?�Oj���3��_���e�,K�y���4���e��h�x�I=�	��K@{*nvt@D��~Ħ�.F���(��n�ѳiڽ���f{�-����T'�vC�`�/�_���"�{�r����݋�2"$ǧ�+9�[������Gw#��H�v�V�"�������Wq���G��[E�7�y3v�6�kswvl��i4���km�����g�ه�,���Z�P���js ]l��Z��B��]\���!��kN��9��K�b��������V�WG߀>�.1]ҘS#��lS�oZ`>���cƒ  �:�b�C�+����]����Tr�#A�-�kN���,����I!��cf/�WB�ˠU2c�O�J~���B~���I���t��x��EZ�Q7X�R�V����~'T������FC�	��������5ڂ1������u���W�]_�=w��a4p�6'��b�<O��uX}��E�P4yZ�g^?��l�+靿5iR�⇫�xbj2�nS�P�e1���.]�0όձYY}i=����䅺&��%Q�����,3�[�:9��,�-�ɉ��D���Z"��^�t�b���$��/N9Z̅�}���e����?�K��,�ӑk��j�:�[����FNh��z��j_$�вO���g��f{�$i��e�K��"U��!��i�sCb�I��>$`�� 3 ��5ެ���H����P�F�b��{I�ї%=:�.�k�L=������N��Aڌ����d��u퇑���R�����3OTA�"�ڰ��c������������M�3��q�/1X�2��P���6������A�t�'NQ���`jL嫚�A����W[5���Bw�j��������=6��D���ǳ'��{���e;��=��rR�\����^��E��p������'}6�i�ٔ5�9������<4�cSZ+f�L�4Xԭm]�A&0H=�D���Ҡs 6I��aWY�	�L`���	7��3-�ۚ�kx�O�?UOP��`�J�ۮR�e�h�AZً����U8NU@�3�i��C�׬�P���`�y�����I�W0&$�I(JH����vS�r��>y>�CKgSl���\��'\�_�ƍ�j�[~:IT7i���1���;�a��j�@��*�ʠo�M�ǎ�r{�,�F_�m�'��K�uR���u�VNm���Q�ڹB�ե�U��d�~�9��t��I�g/QU��Ѭ�0��cmm��#�>/�72��Iۣ�2�r_0�ө2�Wm��+��`�Do+�$�:,x@l+��<wpCxĺ-!k�f�e�'(�����L`��)��	��l	��ә��5��,�Aĥ?~�Ң�Tx=�j����E��}�&C��gvF���}{S�=^��,/��?O���n��L�5e<����3���6�AM�xn׏��?O�,BN�hJ��7�z�B/�3^��Y	p�ȣ�MT+�ߴs�x�i[����sS!�=���p��ʬ�`>\��2��ž�J�/�^S�4ׄS��0��j3E@��aq!�yBڽ��}���oT������h���n��7ɰ��;u8�:��˸x<.nX\8;AP�F�Q܈S�ƪ
�B�����Qz�����PHxN>��~��{��	2=)&T��Bl�&h�Ђ#�F���}���1�S�%�/̪�9�_E��@���w�����Y9Nd�&�x\��~�π忀����w��hy��v��^g�p�19�*�0�q���T4�G�ݞ���1�yނf8ļ����9�f�fK�g��ۉw"n�Ҏ���y�e?$�{]_�J�N2 �F��2��X������:�t�(ٵ�������45$���q*�Z���)�Z�Ìgr�S	P���
�E��K-��_ =y��	TS�����EN��b��Fپ�Q>�{�q�/K�1zeܵw�r�/�l�2`y�H�X^ww�-j8��3�����w�Z��RO����=%g�7�]�o����".�?��H�`���aeP�i�(��A�8�$�>�#��1���H�$`U9)���A�Pr�Wwב���Ze
`�eB�Oe�n�0��U1��>ŝ9����Z��������&7[��`sʧ5hj��z�վp�*��d3��)��xG�'e2#��	��@C�hV���dv�����l������>,H��ֶ-�&w��޵�,��j�]�_p!���0��m�1��f��x����jY\ɏHƖ���Op�vŔB%<zW�YlO��w����\�n����ɧ&���GS��r��|�v�:�ޞ��{,�kZK�7G��vo��#q�n��^q\Ky�Q���seD�Ơƺ�=|��V�����n�`�������sͣ��V��ay.8V(�	��D��_�Tʮ��zɠ�v�$�:�҉70���✫j���8F���u�I�����/"����HZ��x�m��B�������a��I�#<�FZ1Z��!ͫ"���O
�w:��`�9�&^��>�7�z�I�3����v:��8��єN�S��H�г$<��H�YuZ�E~�}k�V�`|�΄J���IUd	R�p�	A`�6e|A7��V�n'z�Md�j)˪�<�!Tq�>J�������c^6%Qqs� ��+mo��at��HP�ѓ�(��~ �P���?�L)�ŰK��2v�(���8����$�?��xP��|s6�e����Z^��-���9 ��c��1Y�1��#U�D���r�,6�_��!�>�E��ū���d��x��y-߻�g燆��P0��GVC��S�q�/�<F$m �&�f�`*к�B�v��n�Y~�c�ՁG�?^�#�pLWD<��l����k�ee/m�6FwgcmTs��L&&-���|�ںX��ŻSXa��\�y�d�x�l{��;�h���Ľ~�_C ���_������q����Ci���B���aDt["��ϧ^S�|�=���c�s��[�1���VZ�e�p�+#B����`�,3)%��X�>C��h�X��²��@������z�AB�U�F��H����m�����O��"��\�Zy��`s6��cT�V�2�WH?o����N�U�4Y��a�K����s�!�s ��+�[��i"���F�kP���I[�I�;��H�ޣ}��1}���֍dy[/§y�7-�Ί @W\a��-�t���PҨZ�"q;6���F�1FL&�hJP�4���3?�N��jΒ�.˨��YIm��bLO(]~-8���KA�?vN4�����M!Lx ��;��lC����������;4�lEMe�#a���l��2�j\(/�l}��U�O�f�'1,���	4A���N}'!�Ym�lЋ7Y�eV-��h��+m��2Q���Ʋ�&����h6�Z��F]sK����VeV/2�O�����,rl�`��ݚiR�Y��^����𼱀�y���ǟi2�+>��X�3 �<��N���dt��X5�����Y���l�z��.���ik�)�y��*G�]����<O7܊~to7�ʅ� �]�,6Ձ[9���,�f��(ጝ8�Ҍ���, [h�N����ՌC��c<:�ݝ���hD������I"񨌽���fAHK����k�mW=~�"+y�twvDQ��I�Z��'����d��LiF�&
R��D�>���1@|�S� �!?��v%�r����'���E�5G��s%_��BP�[ᩨ��˛«��s�l>zE�7��qeE��l��V{"�-o����]ײ��Np�(	><PO�Y�F@܅���/I��U��TS%
���5[�sd!뿪Y�e�Fx�Ćd��ݲ�UfW)F�����>���H��!�����>���wx1ӡw�5�0g|0�W]�p�a�
���+�+cj B�A c�Wox@Y�g�z^�a���2I��[ޙZ��_+�6S2�)���:�E������Dg�#�5�7���{����7D�[��IS. �ȶ�d;;�Pd׾����j��ld3jM擙7M�~\�.��)�
�ƁΊ���&6ܱuϐ�@[��^�����}�V`e1݀f7^,'�}E6�Y�h�*�5�A�@b#N���V�R���?�_��=�Y�G�����P?����1�ֆv��Z��{��%��yM�L{���-Ҥ���~q\	�}Y-cO�;��(��-@/W��ۨb�l�m$9��y�x�{4��u0_�WZzw�����|`>�~�2��6�Q4(/�!��Q7���Cd��p�+���w��%�&	�V^�6��,��p����TJ&%�����~_�W"W����yb�57V� R̖A"@d�T^V_��$�".��p�ge+@��f�K ���'��r+��w[Ή,9��!0Hڗ�m�2w3�G{Y
��~�M��9`j�$ѫ'6���zn&9��hu�5������H6v/�ٟ��N��)c�c���F��J��������0�I'f������zy�ןS��c�$-9M��a|��p�52����W��pķ�"�#C9��y�gVw6��[1�#�B����3x�<�Z?V�_���zC��'�e��d�ϐ��YGO�c��nmÍ�ϳ�p"�N�<��!��[6j7����F6�x>�'p��Ef���9�=�b$���Z	P6��/H�
9�ѐ.��<
��eX�t�ć��	��$�<w"8({C<)�G��?�_�Eu�'K9��Y��A9���2�����nA;��a�?p���#{�ؤl#H�}uJ���@%����p/������*	ǽ�������ԅr��,�~wa��B�k�J��ɇ��)JV�o�*�O���	��u�9$^ص�Bs6�鲃{b��*ގ��K����Y��D/��"�+ZO�
�-zy�*¦���o��:Ҕ��m�O�k�q#�O&>��Χ�	��va�Ҙ�+
���QIh�kg��(�j��D��a`P'���>��f�!�;\����a��s���\�-/u�%�X��6�-�.�$��LÂ�a���U(O�<�eF�J'k
i�G��	$�YF�g2��/pq��R��R/-�[y�����tm������L����#�p����=Fmr�����'�ͳ��[Wvߪ����r�ҵmʍŞ�"c(�;
:7m�F%?�:�jtG� G-�Bep\"�9�^�ȭ�p÷��7Tѐ�)�v �ڢ��8��{D}�ڛFչ��A�e�@�w�Ֆ!G��d�d� �ح揤�S��d0���ã��bWیB���.�1i���Pھ���E��t(�4$ש��:���7�;����b�sC�h|@�g��FD&��1d����_��.Y����+��H�'@�R�7����zS�%݀�tb��i4�V��<U�1�w�x�tg��1t����ׄ��5�c$���n��Q����w𣸀�g2�z��c8�ς�4?(�U�H���9깺,s}�Qc2BY�:�e�{���������z.����.��j`�J�2a���Y�(`X����_���=�?��~�dt=�j���5g�'Pn��]�1s�f�K�y�)U*Jk�����6_yF���{�g�A�͖#..��E
{6�S-��+-"1�p���p'�[��w���\K>ٵ���c���o[��@Aq��#�k���J>N�.�2y���B�pHR6)(o��n����U�����%G�c���~�Xu7�ʺ��˕Ý$��j�RB���t��u�g�(�\8���&e�����00<~����z9Ӎ��B�|꒜��ZPw�3�3�>Qn�Sh�i���cw�P9d&��{�ͤ!�a��)�6���Y��Y^uB�Z����kR{��5�M�b_����/?*~�[G$�(���_>:%�fr���6�S��P��Oλ>����p�l������>d���r�����W��1�fKq��A�y��<�����qN��J�=���7h�z�VxPH���u��ۉ����(!{���nB'#��|(�]��|{�e_4e��:��س�n��#G�܋���,�J�R,�Ǎ�YYIG<<�-��eW�L��t�sE��d�'���+O��C�=�^�F��^ٛ)q�jl@����G��8�b6u�A��+�M�DxR�T1���Ƈ�n���J��yv6�����U수�7wKnˑ�:[LQ�G>���+D��0�c�,�!����ΤŜs9�H͜��Aa���m�pb�=!��"(46�b���mRxrI�ѕ~�?R�O����
L�x��t�I�;�^U�H�\'d��$۵�r�_��cu�kso�v����ڗ��C����c`�`bDrq��w�J���q���cS&]��b�4���3D�Ӑj�|��	_�Q)�΁U�8�TC��E��ǧ�����A *Qją�94y_C��`w5����2=�;��dѢ)�_vyd�����!֓Mi!�Om4�)*>�'yԆ��#>CEh-� ����ke3и|ә�D��� ��3٭��wU㤅�p�V���i�d0�+�����ߏx[�FT1���u�_cH�H�����bq��K@�r�D^�/����܃̂�E��:���f����/e�h~
+��0���o�~qj�DWp�o[=�u�
�
��^���. gp�5!�{��U*��J�����,K�s7�Gt���c��#�j�B*�-�`5+�����ͣ/�n�g�`����jK��h�������[#��n��$dY2����ܓ��}M~������eeȀ�^z��L��ڄ$-J����@ ��C�ug:C�ل�t�ǭdv�
:j��!�K�)�#���}7x���qX#Q"�x4��rB���յ�7h�]����	pV0�X�9b&�qC��^�`U}I{jy�N�V��_���;���&�;���5���1��Ńx�+��#J��"���;��(��1��}V�+f�X�f1����|H$� ^:�����	��>
Ý<�$y�TL�v�n�U�n�T�T^_��(A�5U�i
�8���J�S5���_�������,����l|�dk��>�����W�F���
��Y��E_�}��jS�@���b���O����0Kѵ��3�q�蒬mX��ـM*�+�ų+�,����#
V#�RKTJ������u�x2��@bL���AͻG�cFډ��Gq���a���m����׫E��4�_�ܜ���r�0C��8}�]It��|�^��	�Oq�������dc�ܘ���#��f4����Ϥ'��
#�@��+��i(�
|�p;0��LD.�2I��%|a�u���g1��46s�hƂT�Z{ݵ���p���^ۖ���ũ�NY��6��o�5�C����=�4�Ѹ��`X��)����d���æ�*=esZ3���FS#S@�sx��cz&���f����~В���N�-�\� 4�ҨS3Edk��;vg$��� ����4O׿���IVA#l)\�A֑E^  ������;(H��e�����D��]�|�m3����!r��P~~@�Z�Ci����g�Q�Ϻ�^��g3*�缔���q�����֮�[��L>���S�STn3��:��p4��_�Ly�e�%�3!�ծ�7��N,�Ⰽ�X���~Ň���y�/&�Ha���\��,��O+gf�CEw����c]qW��Q���>�J����q���n���򖯘�遍���.rG[��(����9����as���J�*�;<K�`��8���k�9�^/ҡ��9hPx�]�h�mڙ�߫fs~4΃@�4��B44��ߔ�3��#˲��]	�dH��m,�˱T�é.v��O�5���t��7b�z,>������<+�&Mlr���yv&D��'O��ٷ*�=Ꙧ�:��m�����2�L�_�� \�L@�����,��U�mm�m.�n�,4��P�]o���!�WS���[�����u#)p�R�&�L�F��d�6vxO�u<<YZ}�P���z?ή�8��)y)W�ݚ��