��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�QbQ���'���rcm3-�m-��fڃ~��:zq�e���P�ac^]p/��.�)�b/a&l_�5H�*�k�K�!A�ɝç%\��m|��YY��"E�G����/����+���;�{�j�2�S[��H|�HV�uL��M�6ޣ�R�\F]�E�֣����I����=�N{��5[F_P��/�VO���o�5�Q�%~�]��)KL�L���z�XBr���ظ��r�C9VsP,���j�t��`4�&BPhQ)�ׯ<ֺ��T���/&n�E��$��ۓؿ�����!�jp�H�Xh�*}����I���e���3�̲�q����� 2t��![�>o�U
m{x>��P���?I�$ȫe��w��2�l�������w���I�nq�����bty���07)��`\�ku|�ي�L�8��L��O�%��a�U\xN�f��(�:�6i�E�cWN@�L.D:���Z��C�$[aXД8yw>fׅiN�|s��F���eG]vBN4��]߃�ip�*�ͥt����#�ЃC�i�k��)ьx�x��y/TF���}�xIW]��^��o� B��{R>�0��G�����	��B��l��ў�f� �L�f(ܦ��U+��nb esI�G�3��~_)��%j�)uĵR���E�3�'��n�$�'�2
�.]Q�z���(f*qČ��*=hc�g{�`���{�#]ޑmA�?�� S��W&�䘑��MA�z��$p��<Z$/���32��6��%�[b+�lR�ĉ��B���QZ+���r�};�Km\^��X�]����FÞI�n[�\��ԃъ��O �tϾE�m���ᶠ�Y��4#����k��O^r���M��ɔ��a�)|�dfR�s�����|��h5�9��"��U�so�*���Y�2�'�m@p��H��H��
�.��v�r�'��d��j�ߦb8ti�e�!�a�)�EͲ�E<���ahT�L��u��?4�4��*}���s�i㬴��r_Y�V�ǎ����wW�<,�>e�X���;Q�l&��uJ-m!�_��gg���a,8�G��}J�tMYIS��eW�����+�N���=X��vGpU��-!�v5zM�.�۲	ձ��)�QF�&Զ�!�9��2�B��1k^�W������l\A���)�̲�]4���?�O�~s�>�g�N[�p=�k��$"�û;} ���ؖuUI�Sԇ}h�,˶-&�{�҉�����v.�� ��'@�.��	�`�_4Zc��B�dq��n�o��� r�#�����Z��f�>���&�d��~�U}2��,�ES�,$�r2"`k��9�~'����lY�l����H�SA�և��������SϙK����I�!�z�3��'�ȅ��]��#}6=Q��Ho�g��R�PC�_eKl�cU��%L��]��&OU������F�2%�`���o��ˬ^���x5ޥ�z��.��'e�B�����C�a�&��]N��(�'G��U��Q�.��'x� z�F�"ERS_S�� �P֪7p�"��y���˘5�J �/�U���
{D��}��~e�h�0W7m��r~~-
;�YK{e�=�O�D�z�ʅ�{g>G���Y��b�:4��8�hj&;*c���$��Y�	0�cюA�zsH3��XxS�0բ���s�7P*�lB|&it��Q��U���R|�3��"�rsV��47Q+���zٔ,��;ڍ�����Έ�i�:�~����k"�A5���UT.ORϺ���cD#�ì�:M��tWs7�Wl���w|�C�+���`z�Ⱥ������LQ��,~��P���Y��x�O��������DGtsb�?�p®��l�뙭T)�7 	R���g�|p��qX��i�-�^̑���ë���ṷ5k����'�B���F튦�X�.J3
9I7�>`�c��1��aom/�NÙ��3�P�vB\�X���"���v�z�q	�����O�!������}3I�JNИ����p[k�6�*)!,���ý��B��)҂+�U��c��3]�z3�m{p�A�V�}�3����,��"���g�2�?А�l ����خ�����%�ؾ �l?�W:|Ѝ����-���a�ⱥ�>sLc�E��{-�$j�"� �B������ɞ�>��u��G�������c ��$X'�f��B�Js{_I� ��:s
v�b��Sw���i����z?�l��&6��������QC͢r�Xqއ�l�G�όO�vI��܈�sv�]I�a�mO NS�LW4��3魯A�>h:I-�2Ct�{�GEe�o#��jx���dX��N��wɌڦ�,��U���w�v�1��
dP��]��Dk��O�/��<W�
�����ա���xy�2h\��ȹ�&�.�����V:��%@�GזPbX���5�^�
�\����I�����>���w�7��b��HF�����ט�'�A����fN{��#R:�K�E�@^�α <�A���SJ�(��+�P�,��V{��WA�)�B��;�� hi@vlaF2�C![���"�ҋ^���jc���pl�J7>?��".@���=��V��SM�j9o�o�~%OR/�*�����?B��o�I� ���+#[����``q�,����=q����.�c��:�Ơ��T�!��|�{S�v��'�����f>¯�.J��TM32%�5L�"�J�<T��cz�Y:�#��[X5j���|X��4��Q��v��B*�����ە,5�'Y8lW���zO R������Vi�n�s7)�(��Nw9�������w�޳=��Q&Z9�H݉
��
A�'z;��$#��qPyǦ� ��0ߑ,�wP�XXn�5��W��uut\B$�������gW-x}�`&�+�
���U"j.�p�X��
�0~;0�(��Jb�2@��M��U��.�ӂ?Y���cIn�_~	�p��%�e��y���[Y���ŝg�EQ��	� ��m�'�m���=�3�N-L�[!OG�0)D5·U�֨Or�C��:��<֕��
���A��a��1@jc�=S�^��O��̑�Ya����K���OY�,ۄ�}��Z�{�1��w"�bsF8
�	N�:,�E�͡{�ΰw
�*���,q3@�#�n�!�o!�lHG,�Qd����f_{�O�$�u��y��3#+_a
�qr�l��LSӯw�K���G�P9tڭ��KV�@�Y�
��n���m~���4����b=�|���NB�:1��]�	D)~٨檷�\i]y"����{|7��_W��W��#��j�h�(Ru��+���5�#l�}"���R[;_�0q�_Bx��!��u��a��ў�A���B)m�x�.��K(4̳(����\|�%_m)L0��{sC楣(����Cp·S)C̀�I�#��V/���� �7���T�}�I�i�g��k��9��-IA����a��Rd�|4��\�:��8�D`Dm#�?R@y�Kw����7���k�陒�*���b�anf����2WZ|�r}8�V�{�f|�l~��j�|m�� o��}����%����a��{��y�ð�!7�Ѯ�-7�?B����;���?�3����)�.bE��K)p�k��3z|]�),��a	E���;
��JY��c�X��mו'ON����>��kt�f|j�K�m��o���Y�c��߸c�E5�+4�'݈�*(N=�!8��K�.���� ����_��m3d*��J1͢��7�Vȥ=.�r4�^=�Qφ���:"� �xwa�Fw���Vy�БY|4�>q?�H�N��,�������}�X�
���Q�Ji�'7MnA���W���6B7Z��H1<��eH��;F)��[<ǰ60Z��z�jq���OT$,���¿h:��:�Ŷ�d�P�b����F1kaF��O�S�_�	�T/?s��#��NC�W<�'���M-��æ�k �(��ޚ�����a��5��J	
��_AHR�\D4xx���O
��u����U��L;��l$=@����c����0�p �/��洌�m�{m~�s<q���en�N��_�y���l3DߍYB\�񨳹�a�#I'z@���/�dzu�#� ��:W��(�=��:�2,p��n^��h�!�!5��n�kȄm䬸��X���-5(I�F,����"���"��u�h��?�=��jO`�M,>���._��"�<D�B7&��$��>��-���3�P����r�F��w�Pi~ǣ��u)pq���	g8~'��X��������x���4n(�EI��QsiJ�{k��3�Ir��\�2-��tG�&��Ȣ�>fiX��wW'����I6zs�/���X���C��<���R �#z���w��iK�E��}��2�~oB�����a��W�m�U��pW�3��UΖ\7N�yM�E�ԅd(5�v<9W�+���d���¤�"·T�j��r�u�a:�Mq5��b��>&Mm�=��ӯ�δx%Պ���J �ժf��s�$[��]��N0K�j��U�ʍ#6-\P
}��@�m@UQ�6�5���`p���7�t.���2Dr@qk珝�-�X�����SBD����V�e-4�r�)�U�Ec�8��'x.���	�m
���Tk	���a�e�,�GN����@2�����:cyJc��[T��ħ��*�'�"�8��bbѢl	;\�)��V��_L���r�(1pN� ��\3���>	�jͣ�f�VT
`5]����y�"^�[��)���.��7k�\�G ӊ�^���8�m��ɚ߽��������c���y�%�pVѼ[HB��>q�;�I��~���u��u�M�Z�=�JM����@��L�=���yʎ��b��K�LS�y�Oj}����I罦'���񨾛B&m	�����ZI�g`��[�_Ī���1m�ET��$���7�rK�,�bc��Ѡ���I/٥��_*��Ŧ���d��h}��r.�7.I���i�� �L�+������aJ7����[;ҥ%~�6с�c��W�[�v<��%����"	�{u?
'��V۰�8d8��?p�my�E�'�gT���V�M����Omm�����b�o�\��ź�� 4��Mk7h㩈޺
�A���&�F�2�F��sQ�9)�_�j���o��E�e�kփ��c�!y��Q�b��&�l]����UI�㺽�v�2�������Nj3@:~E�U�{��Pk`i�t�̭���Yh���j�Pf�(�*ӳgNɝ��Ƒ`�KUD�k5��|MH��@Z:�[皴Xc�	<��f���b���a��,�k:9s၌�>��4�Y[&�Rq�RK���%�� ɨ�C�l�Dh|5���N�2�%���rb�P�.] ���8���S����[	{��?l ��w>����u�q�ӳ�R�*�����ڷiE�'s��>M�A6*&m�!����I��eT�M���c2�S���#>�ujo�@e?�C�wN�ᯉ��ЊѬ��EL�\����X��u^�h��-Q��0a�k&��T/��`U��L��MV�@�n�v�ʉf����`}=�V�2'���أ�w3���{I�Lͯ�=��Syb'e"a����*�K�,�,�ʮzy�XӁ+�h����;ůf� ������B(될o�?r��"�Gm�3��:.C킞��j.����[��@�fUW��%��Ժ�~h����Jn�O)���p���5OL��NL���RY��jП:�@��!;�#�N����/��|Eߑ�d�1g�~� ��n�v�Sl=}�So�S[ai1}��s���>�.�2�:-�/�V�)����Y��п��Kj�0��l��GjO�0�yt)��ƭ����b� LH�+5.ʣ�(�T���s0��[��cUF��?aڪxu.ox�W�b�^ۨЄ_"�ɘ"Z%��|�9���	�E��dnΛ���x�
9�z��N�(l|�@�/�$���2��(sQ������/®`og8�LL�w�� ��(+��5of������tT$����ϘMe��g��?�I���n�1VlG�n�@ ~�Bܷ���L�|�!H[�a����y�7���l5��br0���W����N1�dJc^��p�1E�jW��k`]�K�0�8��fi�>�2r��ĕ���x5�<�r���?;��g��e�ҁ;	��M~����-	�ֶ:���������J-�z��ӫ����+��m5G:�&m �2`���0���AbǺ)�&�����$P4�@�#rJ��ojLk���qf	Y ��85�(��N����wu5�*�2i�#&���b��}�U9���4��$�=�_
p�7cؽ򉊶�ß
4D�)�@(x��A8��f�0�k$X9���K\;�<j A@��6~1۵�?��D;�Cn @�S+�왪�yt�^���ҥHS�MR:Ϭ�ւ�h�K""���D�t0_솞y=��D{�0Jd����X��~��Ådd�sU&�Fm��U��rf{�W��YՁ!w�Ε�Y�5�t��X׬��iH���@�P�ʅ��q����uĖ`��*ᄐ�{0[�һ�7��!���K�[8��a��rFRI:	=�呵�A4��{���?����4�2��9��(a�i@:�O�T���<�%��!n=��`�ɨz�z��Xo���^k˻̯#J�z�nЭf��s.2)�J<d��W<:�N���S��1��������m���4��m�t�����������Cy�,��]!�b�Q��ǈ�,Eu�Df2]/7{��kb���T||�s�ai��Y��=y�]�bK���gŠ�ٹ-�� |���8��uŨ ���q?DӰ��p\HiW�V;��߱��!��"��x��I�`�R�Q5r�Sz#a��8$ԝD�"W�1����:��K�� (��ZT����Ԣ�?�Rӽf�{E��\�i�h�f�IlW��k�;��Y<=�+?I�{H<� �Z��#������� �������q6[����7x}��`gH��N�Hj'���!�h{�.�cY�D��ʠ�� g:�'�--K��9�.�HX�9��/w_6����m�Z�_ �='����� ;2\L���b�\n��-��E���E��c�V��6V����;v::��õc,��Vk��-Mv��MCPS��)�1Z��w-���$��qkև�.Yz����@k�<Ҕr���WK�������Ó��z�qޱ�?�i��dFP]��	�΅�_�����7%�|��������u�2x�HAڄ`�܍�Zb�@<X��@B7��`��Z��T����d�sr7�Q'ھB��X�Ue;A`m5G�l���u���1�=����<��א'�Q;*�c�^v"�������Haσw�K|�I8�YI��[|䱧�^#��x?4];œWX�s.`�-޴�	�����$�k��UjŃ�a�X��h��c�n����0� oU�:�xg�K϶xFB{�r��	�%�)�o_W ��AS���
pG�E;%FJ�^}�"��j��p}��]=���
�|��n�-�n�v�\#�G��Z��_q�̅�R"��m1��=��k-�����BXP�0KG�WW����uL������A�����*Xmb��A���P����s��ʍ�Sy�<��KZ[h��_�U�y���2��aƿ���lfޮ��cV꼉K�tH;�!v�A�(��*b�:$%������V�"Pm� :�&���N��E���o'y����4�TQ�
�z�x#�5E�۴���0�{�<��8k�p�y}�ˏ��V���'Z%���r)��Z}ź���,F۞uF�NW(�	u�gI�N�m݂�U$��;BZ2Hbj5����Q/M���xzR�w��4�zi,g�_��w֏���l�Fe;�+�N�_�&_���[1k�k���,O]��{�C���Ɵ���UCf�"�Y@�x��<ƪ����Yn�'������(��[;���������C�����.V�S�vi��&��Q�z���8�~���m�di]h�Y8=�km�OʸY�,[��X	}c��0D�ɏ#u1�3�M�?'���WϦ]��;- �H*_}?<A�P;\Y먈�'V��U�x)���l��`�Y���]��=�p�\d>����|<Ex ۍ��v8"�����)�e��L��fz"��1�(�jAGY*g՘���A`���*�b�
������G|�7��P
떃��x\u5q2�;�����F�	��T��T��]��L��k,w���ܦ|�2��L�O�¨��r3�6^]G�=.����:�l�o��1�K0j�Z�n�����
���=5�z�Lv�hYP�pn�������g]�=S_����b��g!=TϾ��d�~ݘ	e��B����7��Qz@��Љ���Z�PD�Ϳ@&�X1�~�d���r8Y���1��hA�}���O�ki��4�lc(�l����{��@�VȄ�3��I]���y��E��I)�c�B^0�vj����㔇,):��7��H��}����n	4����|BX0���c+�����J��)���Y-96��[��^�/v�[壡ĝ��[۝��r$
P�jg�M0�w�R���)֊�({<�IY-�ꓔ$��~�@��(_e�X�ftNcm 0�^4��L�N�A�*#uյ�s_8��]As?�w]v}����d��d�s��$��҃�y�8u��{�ꄽ~��?�k��	8*;���K��T�/���e�@8y���*��a{ ť 1����m�kk �����W/C�a�����d$�t�2w���#2�<�a��&�J�wC���� S��`d@�j���l�9�̷$@N����QYH�aR���ækL���[����w�i%$�X����vK_mkuˠM�, 1:.���NA��{0�B��8��o�$��!���l�s�g#Xn(?�� �¥ԃz���uz�J�k��"��b6�. ��r�f�w�|��Ry8m>�J��ozኽ�6ҩ�����FZ�z��S̎E��[%��s�LH,X4%-�dCr��I"&�����������:`�)$�e���Z.��A^3co�>g3'S��C�Q��Q� ;���(g��L���p�u��"wĳH���XQhȋ󊡿U���ɑ�R�TL���,�WT3�e��,A��q�����A����*�׬�����9⁛58�2*.�u�B��q1��
8Α���^P����ݻ`�3*Y\���t���}���0� ����iX�%`��	�g�W�eds�F�>������,2=��fҺ��0�[���K~,�A7vv��P�>�<a{	s��a�C	��9b�D1��kKl���IR0��C�G��8H�xK�%p��Q+�	K�8stҎp�S�D��0��+��L�d�O
`������9��zKnc����]P�x'B√�p��S۵�������,�W���GZe�F��/���}{#-J������������dU%���'4�"2�*����v�&!�ʋ� !]<��Ή���ȅ+c��m�ž�� z�?t���	�.�����h�!��Mx�ǜ��ۊ�`��I�0X&0�yh>HO8a9���>��a7㙅"w���ߟ�@�D�����?���Qa�-I�9���Gʇ=���)SS�k�Vj�|���_f;G0�Ӳ��2K�ns�����Sv�yl���(*��r����6��si]w���&�3�}evZ>~")G1݅�DoB�lC?^˾��o�BsC�"M���4U�����Ty��Y:9_\�������@��N͘�F�sa��`)60��C~��ɓ<�yJ>|#�cc�$N�.�v�};��dH���0�]��}��7��R�o�N2+1�H<T���43q�Ϟ�&,y�w騺A�&�ft����(tX�k������T)j#�Mdܗ2��R�Z���؁anG��:$��Y�a��8����!f{.X������	^Y`b!�C1�gzx�r���mw��U6Ah��]Ҿ�C��ּn��V�N
)���I�������ݹ��e6\��L��S��z�:-b�қw[7�"d
�ᗧwU�M1ޟ�F���r���8���+5�Y`�}��S��Q��=�'�Ǳn_|��-�:������c0p|�" /M��u��6�U���U(�s /��NRw�nj����Y�@/��>�Quf'$�
�T��2fى���޼��+�� l�m��G'�����$b#mB�K�J��]q�+����_ dO��\�87�Y�U�����
��^,z�K�>/���|ɋ=�*���"����ta[��&�{I)�%�8Ӗ;��
6�ͳ�ץ�c�V�>��l���y|��C3�J7Xq���%���x\���Ofx�͈90��)W(���!� �;�[~S�Q]MKW��1'O[T!�ſ�`����K�
��܌'�P�-瀨�]�OW��t�T�dWp@��9�Ǫ�棎��nAA]2��q"3����S[C��͍vbٕ�y�S�8Y�\�-��i���Gφ��5�� �Z��s������ }2+.�3�#�[�k
8�7�Je�ڑ�]G��e~n��T���)�M��ZlAzi��_S{x�X����*?�ni�r�}�a� 	8���&����hxhԤ���=�n�A�R
�:��m�d�G?��[��"/���*1Lj��	U�ǃ_���.?f�Q�<U�3�}8C��Nh�	߄�^�j�CFr$��c,�>�QQ�}�H�!)S���>%^����}�1=Q�.�y'��6 ��`Y=g�ܐ�T l�m�%_*���@����$0�x���ej�y��?�:���	�պа}r��-9k
��؀���0I�h:��2J�D" �ضN��$z$�s�M��@�r��@���U�)�����_U�0�Y:��x_��!��'�$���N����D��Gkft��?�.�� �;3,�Y��%b����;�FT�Ɏ���ļ��`J�&����0��)�q������䜅A'��X��Q��<�ŴW�� �I��s���k,��/H��Ρ˟��W`7@��	5���+դ���١-��e�0�8�	�'�\�l������	�%���,k�逴�ak��%�U�X	���-]K�Ͱ sY�bz��C���9�ᆽ��9����Y1���i�����K���XubM���G�B�J5N}4��W���
5Ӵכ��y5?eQjd�'�?��h����k� EX��$Kg�w.��r���r.��j�y��iI�`$�ǘK��2���~w����ju��ީ��[�����OQ�IcҘ*���ά^�Yff��&���B�=P�R��Z�G����Vr�=1x<��3�S }@LifY���u����E�	9F� 4�"�K��Λ)@=�4�|=@Ib��e�)�}i�|�Cٞ�\8ʴ��g�}q��Yd��&(��[?{gI��b$n��J[p��:.R�� L>�?M��/�AJ�LW����S��>��|�� :Rt�UB�t{n��cDK��֙7G3!*r7�ᯋƖ1z4;�v��%X����b@���:��$�Z\W��� ����6ǌ�ݼ�qs�kӑ�A�%�I�RJ:.xۍY�XZ�\��ȕQu��-ز-����,���B�{Z�p�8!'1��Q�+%��t�EN%�1�Ƿ��3���Ey^�A�r��.롰H��L0��b,�
�)��s���y����r*�;�!�����=Cn�K�K��V���4�>
5򑀵�cˋUkJ3r�hWTWϡ���=�^,�e��91Ǧ�K�$����G^& ���� � �[0�>2��%G�*��y}Re�j� ě�!b,�:^*F��8io���ˋy����Ǻ�NO��lf#��630���E��8P��(ک�{٧�|Q���ځZ���]��?,��!����(8!`|?e�|�YMV��dU"�1�(��߽��[��B˧t`9��C���ڪm�$Բޓ0Rw�ԙP�h<މ���d��Ē�]�jFbd'9e�-N"բ���0��=֔�u+�D{�	"�eֽ6ȣ��$�B��́����b���Zى��Mn���M ���E���q���;.m�ͭ��(Y�?#��K�0��~"���;^!���	��{��p�D���&.��.��E�V�GB����'���BI�m�k����Aj��&�`Q	��`	z{�;/f�h)WK�㍌��L�~(���ݪ��$<�4��	�M��
������p��ĔWq��+�������u��ƪ0-�L��<k9�g�9��"!m�ED,_(}�l��V����=�y�捋���_��{G&�[(y8����?���ܨY�T� �����t8(Ibr�%�1D`�<���C�X��Bڸ#��yT�Y F�b�3v���c<O�ё1�ј�B��9�sj�צ�K��Ρh�e���^ N�H�݅릘X���R��Cv�#�P��/ap�o�M��`��X]�EJr��תQG�9�Z�m�]��|4���t�Y$�QNoKJ]ND��v�a��o�]ͭ���ڊ.^%�5��V�>D.?��)�����N�O*�%e��Rh�]�2����!����@�L���H�*zY�:i�_�)x�ݿ1�N����k,yn\���.��9��c���X߫۸	���H���⢙�����A)2�r�1��a+YyQ0x�Qj2@W.^�@>}��C�����@}��=/���ʽ]��]r��ķ;$ �1���Y�3��q�t]H�Lc{�Њ�q�?�vN��r-�^B��X޹t$���������Ա��I����ދ��4��T��	M�q�ܤ4��3������,/��	c���k=�-"g�$/���&�Khsqx(�Y��sw�� ��<z�{�˒��l�y���t{��q�٠��`�)�~=!͓l��qj�)X��"m��Z�})�|5v_[��ۻ��SG�9-���肩~t>DW�e�=z�Q�s��m���M�Z��A�A�HT�n[ɸ��ͤ+�i�G�眀>���LD6︝`Z�sЫʗ��q��<�����_�|�ǟV�u��3G�X��o�RV\�����|�ڄ�N(�8�,=�-��l�����;�U`f\�7�'ޑj�oօ�!��4Ǆ����%ʯ��<s�_��!\���c���!�/1藳y�u���g���`"g�w�+���)�T�	yX!N#���L��}{���\��ZaS���3��q;FB`j��2�\������d���.�����	��CM����=�( zǋ�-�/�Xp��-vC��d�Wșѭx����yE2�Z[t&ON'W_:$N�~t��v}��l�k��ǡ�|DbAF�_c�ӝK�
�|އv�D���Q���W8IQ���L���Rn9�{G�f�f���A&��wv�"KO4l���١L^7�2�/���X��6s~�q�X�9`̙י�cHP��>�8r����:s����7�7nw�}wx��&�5�2=��j��LA���λ*��܁4�� �1�����1��c�/#94��i	�b�⿂< 7�H���7aP�kU7-�p��CeN�Vg.LU+�y�$������&.�d����4����A��+.7�Ⱦ�	�Yq�����qd��𺺨[�Q@���q�f+���D��	!�KO������,�Ԑ)�����0���.�D�8	9T)-�Vӌ��'��C�0I��KT_�6��<�����y��t"Ʌ4NC׮��:��WIDb>E� 4��Z�������YW�L����f"�-#�tc� *��3%O׸�
>���:�8����?֥�5��D�5VJ��}�|�( R��@�K�qy7�K|�-~���K�����cfv�-�4��~t�OV1��ϊ�P^�sͲ��ilw���~��*Պ5�k��˜ְ婷�>�	usp �4���U�v�Q�c-��ЅĚy���詏_sl����=�N֎v�oj�n��{��������`d9�s�3��i�)
��]+��R��K�ӓ�[��؁5���cXN�y���[�_���jHPR�i�T��)��vemV�t�y��t0�D��a�l3=}��`�0q���5�ˮ5}�U��v�1)3b�]L��VL+A$ �n�6���;EZ�oƸ�ܵ�,ݸ��vmO�u1qx�ظ�uk�����d/�k�Q�L?K����Omsҗ�'�s~_!8�_^n��mk�^�:��XqOl"�������Qzm�AMf����u�͘��n��N���#���|�/��F��B	����ie�oމN�9�|�V��L0L�N�|��y��8�?���-nLדꉿ��%��ȹ�߻����|����F�H��2X�X�?�mW�A��5׃f�w��tS�G�f�	I��`��\k98q+Y~ܹ*���
=�ɂ�o�w��]-�������L��e��#}�Ah��b6�A��t������=A)��j�}�h��D�3��ԃ��?cE��,�����y
H��g����"��D�ʟ,-cЀ�ɚ��A�V��Ul[)��v�$,1Z���d���Lc���r>ٛ��������s�:v�r�|�Ͽ��X{���:���H��� |||m:��y�o,�v�+���0�3V���Ҟ{�����ޒ.j�Kg`P>o���M*~���L�)�����
�9����݇]rV@�~��Æ�jZN��ߡ8߮�%̼�&nZ�T�t� Z��߾$�-@�'�h�#l���|����B�yֈh��Y�
O��Ms�7,_�̴�l6!��� ����rxSmb��_j�峇���3��t<�m$Zas�d0��re�(����,*?��U�1X����S{���
�9�Z{e0���_He�$>��L����/��ΐ���Y�O�7���"(=!��*Q���-���'�L�r��,D�� ��@9030Ԏa/H�-����%)
�3)�{ba� �1�a�H�9 x�n�'�	D�%p (�+8:�`�29����}oR�������Z��dt:z�|\�k�#V�CeO���$�Ү^G����C��?񉗯K���w|��bQ��C����D����B]�'��;g_�� HG_��P�K��?F���o�<Sp��W1�
:¿}A�l�:|��CLM����.��7ԫ
�t��`#J�[Z������%z#�㜸�(h�J+p��Q��DI�F<�"��=ޖ+\s��c'����Q�<L��	����/��g�|%]�iƢ�,�{*?h;
�<�Yj�*�R<��OR��+�\1d4#]E���0I<�!�� �<v��q����{!����J�������v!]~�M#v,nB��V�e�(��c%�}�������C�a���ǆks�rcX)�j5����w3�@Wψ��ǻ��޴sk��Hoi�l��:�P$]�M4���	���G$���X�_i/2M4�����/Q��D�"S� ����+�.��p�f�#Cf~.�?7��_i�5�)�G�͈`�?�I6�}��}%dG�`�����q��T�]ܲ�K�b]��kn_�c�|�ޭ65A}�icXo�ϫ|1��}����fj�.�S��f�
��gQ+I�l�8����S<�K��q��u��!�TB
<�<�Ʃ��� �l�>��_��S�� �5������xr�U�pr�	�\�ވ�.�%? [W-�NXX�Rg�v��ʭ� =6�z��{�
���˖��̀�1Ҝ��7c�d�d���7|��=�b�uX1MeI����Hn#���k��.ب���-��q�g$0-,Q���9�� ��#����R��HmJ�Xo���(������ű9�?��aX�Ӈ���4y-+TY��.���&��'Н��;�H�����7�<��B�,(�M���?{�=�%Q�7íq���? �$=�����#�Ć��Dր����M4�0+S��u��|ʕdbY}'�2�F�����P�+]��Q�n�Q�%�0}�oS��kڌ��+�z�ۯ��~>�#�7�J5���	����$r(fxl�v�,� �B�TR�Y�܏O�Ǻ�0���\`��"K>��/�\ ~ߴ��V�<�V��'}�ɣ��5a��y>ۡ�C	��朖Ҁw�6(�4<6<�	���
����'�-��H6uW��T���w�L9]��<	=�k�*�+��I_�*�/����]5�	�/�ϻ��^܉���$�G6֛��ʙ9tP��V��u��������@�OR�0uR�j�=W� ';�!F��*��ԯ�'
'���r�I��`��%F;'3*�h�̓�Js#��ӷ�z�>C4��.'����j��ŀ z��馠��<�>Ǧ��"�g1�&$�|
�8�Mb�/*͓�i��c��(0[=fx�ϴ��O8����I�cR�:�s�G��w�J�Y�G��úSd#�@�oEz������Y�<71�!?����Si/2�-�=�@�a!�|UOVV+m�)H�o���-p ��R/��N|Q
Ԡ��7$���/�N�\�i�H�@�t|�5��ͲG�n�p(�is�`PU��3������~Q	�#F]��[½|Cc�Tư��c��SY����o-�I/�
;*���p�(h�X��P�]}���ǖ�0p��91(����!�m�=��3�Q����N��J�P��-�ӗ���ʺp��+�V0�6��^v�W_ W��V�(�SW&w�8y�4��'����|f���:���7�2�[cľ9@^T`��'*���v�ލ>8���7�A|9�X~��#��s�������8Y@Q�إ��w�Cr��A:��X{�虻\�8��yP3��~	,��*�T��:��\�w��c10�Ffץ�P ����	s��%W�8�7"��Q�"����:e7����x؃���p�|yx���I_�yD�C����-r��i�+)\ny�����z�_
g�b�a�:T+իC�=Ʃ���`�8"zz-����ԑ��Tn຤�M�Qp�dV�.&_�$1f�g90A5ھ�d ܤ<l�,�C�F�[\b�v���8�L�+�Ɯ�-�XI�n:��az�1�8aQ#u*Bl0�*�'[�/�f���nnVtF�\�5)�r�`��\�����E�N�2"�	�w?�`�;�jR�'m��a�E���e!լ/��/J8��)�G� �P�q���')��[��%�kD����ࡩ�/� �2"�4
,z���&�~x �,Q!=x���w�������2���{����K�;�;���D�xP}�x��$��ңxtG��Y�[�DQ�S�p�p<���H�0no�tPt{�.�ֹ8����1�J�()}�!��!����]���V~Z�:��L�Ǭ,� �
J����x�>�C�-�����)�'���D���6��ŭX�I�L;��.��V��[׼���v����1�G}%7Ŀ�;�	gR�ί�]P���I�L2���H�L��e�d��i�v 2���y�E`=BS5y�����(c��ZuBL�MTgg�RbCw��w��
�A�b�}r'��� ���&� n�M�EW�z��l,?�I9�:�G��ǯ������^��8�'������Q���F��a�dͻ���[�:�j���X.؝n��ϔ³+��xõ"�|���{L:�NF�6*ǒ�LNLw�9W�`��^��@ĵMޖ�{�kl��oZ철�_y�hG��sxT�
�l,��Hh-i��;s3��K��kIp:���( i���# �#q�b��V��F���&���1 ט��,!=<�x���R������+5���K����8��f����� e�9��*Ԓ�&�����T���ߓ���J���*��.������N�T��k\���ߚ�d�&
�C�|R��8��jnH�V��˭��lKp1����c^���y%�����x��H�& � c�7ܠf�{������U���f�Ё�x_^c	�������\wL
co9���_���=7Θ� �&������q�F�������VB��(��w7���y�°Q�jÿ@t�Ģ��Ԥm�m���B8��`�>0�:�$ُ�G�C�3+%��9jV��^����6�r�#64dÄ����j�lHtP����t{�>G�j���lϠ~�����赫�!x�WHS��J���y��*]�`�q�c��Ȧq3{�U��Qi��:���U�_� ��{������Gch��V+4�9���8�ͼߌ��
y��Ow�F���aV.��(�c�~�.G�ԟ�d#�!���J�%�G1Z�8U�SGj7v5wD�_8�V�ϊ��m�����v^>r�8N���$�*F��,z�<=�-V�PbG=��R�5n1	��˔9k]�t�M�I�|o%��6~�����$�Z$�+{L�l"�|�6B~m2f����4ӇDHpm���y���I�bƔd�C��A4'Ne�������)C�x�R��� 3P��#���É~�1�4�ME^��Ǖ�#'�2ۻ�u� ��%9�g�D�7�H�W�>�f�͌S町d;b	I�f�!:�O��,9L�X��X�{�<�zh�����R��pBi�UQ����cxx�3p��/U ҅���i��D�h��S��FR2,�������;���7�����;G��s!�/*��$Dvg�Y�w���)>��X�����c2،q����7�tr�F���oz!��Wt�B3�z����[��E�Ҋh!b�.�^�m�*�5�5~���e�ii�X���a��l��^�h���j$��M>^��6Y�����:�0ݿg��l���;�:f+4��H����c� K�7>�o"S�w��+{%$b��je~;��<@
� ��f��Ӆ��v_��c��w���`,���6���ǡ,��lX�n��6���[Ii�+.�������f!�GF�4�`Z�i�|�RLe���}X~����9�~+�]�9��U��O��C���a�
�k%O���\F��"���uO��i�?�grZ?]��+"MJc�jGn����=�6���#]0y�n��,�}�v	0��j^�֦��;��Ad���B 8�J�	Z�����a�i��=@�

�
ɽ���o.�� �)é�K�3^�+�{&nn3��_�VFݧ)K��t����1��n�*��X߲����D-�0E��$V̉�Oo�'�E9��	@�v"Pi�l�LA3�O+��j݆�y�J0�Y�ۧu9+֠�"j�m#��;S����Qv~�J�����oc<r��v�*ROs6���JҵB���p��hP�������&c���*"��Ҭ��B)����l<�ڗz�k�bcX�m~����?������@�C0����p='X�V回��׻k���L�e�J�D�Eoqk>�I3dz>y�[����KW:d_"�.C^����ҝ���z8~�����c8��Zb����)��5�o��\���~}��`�,II��GT�*�O��A�}^Ư�"�,d&X�q��8oVv�Yt�2����4�i2_���֠��Pb?�_zOf�Z��q��Zc<��{��Af�R'��O����k�Q�{�E֥Q:N,r�@���9�-�>ɬ����G,Ju鸅�1��PY��-��˿��U ����	R�@�V���FN`���^�.��q�� D���f�,�J?�� Ӈp��Z�!|�`�Z�w^|g���f�e��A�z#sm+��M�g���B�.�W�b�	G�U�Xd��v�����f�z��ךq4�y����'��W:�vIغ
9 !�J�]�;��mHoC��&B�*`�\���y6��Z?���\5O�(�Ql@���!�UT�@�Z�� {9��X�,�aQ�qQ����nL���)�Q�z��`6�ˎ�Rm<�u�<�?u�;y�P�AHn.(��pv��߳a(	ư�G;��	 ��2bp�J�cY#�iZ��bG>qK�ݬ��Es�{9�~��)7�%�O����4��{��_�s�Sn�p�[��9�u~\Z4T��S�&����#��ȋW�O�S����	�����13��N��A��5�E��xXy�*$H�C�r(O��?M��%��'�ٸt�`�Iu��f����n���Gp��|��g�5q�sbrxO��ۅ�	M�-=x�IZ"�b�c�JU�U���̰Ulo>{~?�����V`��E��>��%�Ɔ�g�&8�^Zb��~L���P	�cJ�\�En��Y��u�U-���d䥹�
���ڭ��4��Ĕ(�%2��%�U�-��T$Ӥ��R��-��C?0-d�-u��K�|=>�@|��U��s��Z��ĥ��gՅ�'d�q�`d�Sp��Y���W��r'|h�˜��yOljF�QL�Fq{5�Pa�W�^)S�2��k��</3�TҙPC`Q��F��&؎X���+}_�$�&D[�5��Y8,c�W���L�	A��f�+�ذ�$�d���`d
h���%~�n�/�����Ev	��~�Z`��l/kN �y�h�1�Tw��l�8��|��s�Ny�G��pFb���Y�o�;D<������ٕ��ZK��׃\:�����m�F<���+�r4^��J��l�D�gwx��<	`n���`�K/`!%`q���b���R��u�l�􀬍1��~�_ ����U���bp1���f3��Ŧ�.��\.��A����f�p�ا�Q�O��/�#�jF��W��4�4��oeَ}9;�����vO���P�g�i����EȑC��]V[�ʎ���y���[��K���wl"��^2���BD��ȉdn�� ��u[�H-؏�����C�L����́6��^��@i!fv�LO�G�dK����6��ӉP�t)���oi�3r�̽iC����Z	���+���5�.ЕC�^,]�H�Na���m�p���#���"��]��1���uNP����,�.8 �)�_}�Q�i��)���N���r�ζX�+��>5�,�j����@�U�4g����k�ŹV!3Ey�����'�Sj֣� :]�ހy��$������U�2�<~�3��}/B�"�UN2v��t2�M���A�
ab����qr���i?�UK��r{^���=��3�]�B���%C����E6��Z��YP������x�y��/ŷ�i'оjqbےʫޅ��h{���Z�Ӆ������F����'�⢉��F��r1i�j��^h�v�������/�I�(��p��j�T�Ǖ�HN��wyI~@�)i�
�:`�^�7f0�h� ~td�ʜ��Ѩ�0��>�jyS�mF13�e׿_���k����̥Ψ��n)��L�(��:B�C��!Vm-�V!��\U��嗜|j9��aa���?<�#�R~ỿ���Xg������.v��IaJ�͌�v��m&4�:�8Ѳ"���7�@���ĉ�q�A4������Z0Ưy�務Ȗt�G���2	��3���\��$M��SΥָ�1=���H�;?@�M�X��1+г�7C<�X��H1����|���k����1'\i6/����&a�]��W�=-�(��7�j���[8O^4�v4�Jݺ�k�T�n��H��^�7B��Q���*�=V̦�7Jr�Ѻ$I�T�]ػK�W����1�����7�m�v����r*ܙ'���^���y}/�F����6�4,�@Tk�t�RP���r.���L0�W[LXj�v]�[����i}�六��5����� #�E��|��iz(��� �i$�4��Mw��י�D�.���y��q�����1�9'>�n��-ܤ����_Dl[<�W���_OvdC��:�Ҿu�Q}��l�I�4Ó�R�0�a��b�戳�0��z]k�Ăs`�i_7�1�I�T����{�7��d:�&S��U�������S�Q��l�dԘ
y��	!#�e��e>�ل��
��/���x�
)�ŨF*�>�h�ǯ��
4F�V��EP8�`��l��'K�S�F��#D���6lt\�E�6�Bv�d�;TIA����ĵF����i���[�Mi�;�;���^�"�ހ.H�g�N��?�M��3ȭ���T��k��H^�����h7�q�,�M�0D:��=�z 1����{�d��u���.6����x�s2Y
�����6(�C��T�t=�����u���ކ���#:��,�Ȏ��?[�n���B���X�4��M�:�;�j�y�E�?��J�۽�m��٭u6?��K�_q[�!���
�'��i4o���z?�o<>��Y�~��t��+}�8r�#�2q|5������δ�a����d��EK!���tts�[o���}������T��@�7���B�7�������.>j�%Xi0�z)���>�0��k�t�]���?/��!W��[3=�%w�|"���@XxfZK��2���L
�{����Ct�J�ۑ��������ɰ�-�ʩ�;��!���q#^q�{Jt����]U�S�.����Qh��d�Cs$�9i��a�*-��e�,��`�'��tgT�l�����^�	����\:ڡU�X3M`�חPMih���O�z����0�Es�v��>�]W��jj�t�v�NV�s�,t윗��]�w/ �&�Y�r��ԣ��2���7������\�m�c���y5��D7�"���U���_8=��d�<�ˢ|He`但���y;p�t�I����h��?uPΨp�e��40��ڜ�X��5����Ռy�� c����]~�*Pb�w�2��q�6�LUN2�����v7+ aD����Y��'cjSH�����J�-&��uj2�� �9yO��I� �ؑn�;Na���ϳ<���.�-��l���V�M�-�L#�Ժ��� �c$��A�M�� Z��F4ymc�YO����'�����ɹ܀<�Oy�5�=v1��Ɋu�O.�F/bT�^��A�g����,cM�>��KV�+�8���8��R8�v�>��>�o��'�i���.��6��^���^�U�*6��f��n.մ1���`kׇ���~�!�[ud���M�ꑕ���T�@q����^����t$�NH�٣�V�<�PX���)�Ez�b�_��ЃR��^\~/����u�6Ƒ�������n���D�!��D�������YѫN��D�[��:O�Ajm��~������=y"����h�0��~`���SS�q��Då�#����L�̍��T���B�uj[���C���o���٩���NX@*da�Kݢ�o�$	�=��2-b,�T��|�v���S�6d~Q5�i���)��� l��X��N:���\����4����/�\+/.��Z��1P��*��t���'Х��LA(k��6Z���� �wQ��</�th�[!lL ��M��ʥ�p�F���>E:��ȥ$����`�C,�Yn(��ן�+�Y��T^djI�_�pN@#a�S�b⧓͝x��)n�2#������AE�$]�OOs�ؽ] u�tV6�crQO����p-U���~��{|�rѡ���y���.痚,X`�ohiіNp#H����do/������- Q�QО���8�I�[B�����B���B�k�6i2���b
D��^d���̒	 ij3*Đ\R;������B���������b�A}���o�Ҵ��%�`�G|~������ڿ�ՠ�.�_]a-��j��W�I�ek�k�M������h��_�fPO11�������x�a�q�MR�.Cل=W�AQ���Y�x�)]��m}*Ww�C�@��c�
<����1�:�!q;� ^�ą������g��k�4ʽ=9�"<5��v�;!��ZG�,U��w.e%��ASD�X`�E67'"c�_؋�AN貽�G�k�^]'dn�%����S�m�w]������Ћm׆PE���{_r*��@Ws:�b�6YA�G��:X��K.�!,��<�r�1r[
GY��ˢu��y�5=������z�A��%M�V\l
f�:�nS��l@˸'2��������{Yُɻ�Ơ�˾�R���|���x�1���(�v31�az�p��$6��G�d���}y�Xu$N f�53���l/�C�un�mH$�iI�[e�\X����oڛR@�/�C���+�h�w.(Ώgrx��?�5�&b3H=�nm��(����7L���^K�Ȯ�F���*�X:Z?��s��=��ؚh�uS��t�(��' ����~� �����|�O��4_1K��&� ���^7��"/����/�C�0�ڀ>"̸�\*��x��e��m�=��ov���H𽱋�F�
��6�^�i��U��P& E�&��,\[��:��R t�~�*9��O���$P�y�lE��iL��վ6�/��c�v�~Jr�	($B���ʳ��޾G�~����;�V���ȕ��D ۱�zv0�Uo�M�x'�B2����Fȯl��„ǫ�t j8�r�N��\ǰ����x#���ywl��G��u� �d�� �U��^�RX�/�;���{���-?��{��<A�H�x�þ��� �75:�;}�W�3�q���!�P"��"��arTP�i��t��7,�����H-6@�ߦX�-j���Ո�z�/e!���]٪-id�t�Z��?�L*C ��`������LM7VMK֗�L5��=��|#k��z�x���נ�*c(����b�����T#R�3�	��U�h�3�CT)Du��RO�v�X74q��ר��2����Do������1K����b3�{��`�[���8�F���|��-�a�����²
�ȱ-��|&��
ޢ�YF��`:p�@�[rx}������8�K}�/W�?����CLb��!.�99�Oo����� �;Nr5��M	�Î4���;[��$x����Q�������j؄�x����Ĝ����_�N�8Qz��:���{l�z��wLqg�k�|N��D_��"-�UǰŮ�H0F
+�Y�Y�Imuǖ�Xl�����m������Y#k��pF[��{
�<B7�v|+(ܭ�[c�O�֏�����բ ��?F^���\�����T�Z�G����q<�v@�u��h�/��Ήh7���F�'X�sM�B4�Tޑ�����YogH|�ε��5�4�֙��H1�ӓ �`����l���D��@���&<�Q���'Pf�'ybF|�٢C�ǔ�.���B �,P��Vd��C�{�V��|y��ٞ�Ywv	�#�B!:�[mq�0q=��z��c< t��Ip�:N���,}�F8����_hA���U�v�T�Օ�?��#|@-N�.峄�Q����A�҆��� �Ȇ�۪r��Ӯe=F�4u�J��<0{�d	=��E9�jd��K���#Ԃ��fă��q�g��X_Jvە��q�Hæ-k+7�TwxL�4�G0���B�m�{
bY�4��`Nr>N6W�+<j��o۵�*b���q�B�> _G��o�>4\~bЪ�����L-�����ks?
ĵ�')q�?]�����;|���@�}�'�����Y˻V��G� 4�_��X�����$n$�A��{���](�O��2�຾�w�Ľ4��q��!���{�udɎ��0��K6�R� 0.�����6aD��7:�#�{<�{r?�8��9�]����BS�S��z��{��t����_���<��0�wUy�?���5�f �{v�:$�v��G>�,(�_6�d?V�#l�<#��VY�J�y���K�	z�Xܿ��kB�K�����-.}��A������t��R�7�]xZmW�9j���=LM`̲�G  ��E�$8�ѭ)��s�+���d���e	Jbĺ�`����\QA��f@����g�/>F�'�&��`Y��hWr�~tl`]�n��_J��A�m
����
a��0F%tN:v��:%�?�~Pj��ϖ&$�Y���#,�0�c�Á�Wߗ�X��,h���	3���97Z*Wza��`{
�[����z�g�E8G�����Mœ����F���������m�`/�x�ӂ�����>u;G�Q���ҁ`�ɘGè\A�b��f��a�Z�(�.*���Z�F<���������;�7~K�u���N&(��;֔cGAs�F��ΉJ����^���:��&MS]𹦙��
�hm矅ْk1�}3klN�(���T��EC4y^%@r���4����XΛ�X��e�#�&>t"�hW$3a���������X�Q��B!hyH�T���:�7ҭd��j)OC�,O�[Ơ	��m(��7�����dև�_�Ò��[8ߚ!������������H�&�p��P�~S����R[�����z�;׸`��$�%��?z�]cր��@�✡��U�Q ��ĝO>ι|���ol�ő9ua��΂S�5�9� ��d��	�~jT���l}���#_`�lύY���F�� y8ǰ~���O�8�Z���G��մ�=�N��G)��Z �Wdd��2�l Xɰ`�.��cNf�
^ˆ �'y�k���C5�q&O�A����7�s�5
_83٢%�-�7;�D�|�	�0y�Q/��>��)�T�Qww�����%�&O��.G�s�/J�_�\W�����8��oG�|eh#l3��'\��;�t�����Tu�y#��4��4�%O,u�VM�?��21m�Z�>���X ��g��J��_���"��E������
�͏��������i�|�(Y�5~�9���<�3��*L	<���?��. �_Z��*g����&��@��ƻ;���$�#y��(�������/��P�&2'�D��TS�D�E��7�Z*n��{� �x%��/  ��9����P�nei�1��Cu�)���V��f�`�Ɵ��r+�hya05��_eK{�Ǘ�����@�C����>�!Քr��󴖛L��U�ud�i-�p�gܑC?�+�A��Z�h�\�N��)�N�X����`��eS�pL�	S߈�-��<[�Q��<`ׂ�-*�9�D��g�bEN�x�XU�Z	��=�!?��&���C�x�� PwF�YN����=+�9e��XD|��H�8�hPq��������r��<ܸ6	�1Y7�����L_����e�@y��4���DH�q����I/��&h8�y�$�����/"�YB,OU�4S�8����\�6��T�L�0�?w��x�[kEY�����l� 	lC�sAZ"|��%������}3b�9�*G���)�iF(�C/��0��O��<y�[��݇|�Td�d����7���a��@IX7���+�06�d�xS��j@@1���:�ж�����G�k��Òa;fξ�MB*-G\q�W���`��bZM�	��~ѬE�`FLJ�����'y�l@oe��"XX�h��>�)���qu=��JMH��xp�j��AگN���V-B��İ���"r�b������\w  b{�Ydi%X!)������<J�����'���-��D�J5�����t_;6m$������.���|�Q�:�j�c�=!Z����]8o�͆㷮�A�sŗ�N:�d���E��!_*�H��w�� Kl��/-���P8/z�؟"3z�{�k7�#+�;��r�|@Ҿ�w'PL�'��Y�����Q ����/h@,�:lu�5�@n�IX��@[��mP�m�����r�uM|8�1�G>5Z�W���=���V�d��\[���I�p'q��3T����:�A*�qp��=Cp�
�j�#s`p��$&�]2ڳ
�@���,��+�B�+�7�	#0��C�cN���6��DF����[��A,����$�\?v^Qi��&m��4�	x\����h���~��.�O'�Q��j`Z2y�|DcmN�3�����U;��5�ɗI�PPC����H/���Y#�:��HG���kb8�=|~��ӧ�4����H�52͌U�hi�T&u2@%j�� k����]b~#�'M�Y�o�B���<ٕ�mO���Lُк�&���k�j��ޱ�(c��+&�u�p��f����E�_����ۃW�[�GY9�0������@'ў���'�(��h땞�`��p��O�N܄�OZn�G&���߄<]'?T�(�~*�����*
/��D��]�S?:�*�{R��~ l�zl�IT;��د�6���ʯ����;��1k�hm�����)8[�=,s;МG��
Z�1)[���V�Vu�/ᶐ�e�@~�E��F�u��;Ƒ��VȒm؁�4�:�
�-D����!��W��fjmF|/IK�R�$�,U2T�+�gk(,}Y�4$�F1�MA{ے���t��-�8��.;1X�iUV��#�O*?ԅ�CgC�˔�p�� ?���1U����ݴ�D���Y"�?��Ω���CLj�m��&��>l�CҼA˯{^~�G�Hርח��I������ubT�9��|���0����<w�4'�����L�3��p�yD֯ƈ���1�p�cj����Gq�̋:
}Âi���H���?����Omm�*�cӸl�31�5��
���01>2J^6����+y8(:��Н��3�o�5�
��I�h�Q]��Տ��U��6�,�����"��^l ,�es�a|�.�vA��0�Qʒ6$�ՓO�o{Z{��+2�j}'�=��!�j$2�ҥnpK�Y/��.dxĥo1�=���W}��n���o�|G�K; p��]
W��"���hc��*=o���)��~ŝ-����{�yƝ����r�`�G0�O��(ߚ����6�:$&���Ŀ���:A�w��8
@ј(2J���:����Z��#N���F�]5sҦ��XQ ����)�v|��<��L�1�(��y���[𠖺0'q��A�𣑟`�VNkk��}�p�՛��⪲;4CL% P��	��l�`�y�|�L��]��UxjPd|���b�h�ǁ�N��R��˞���&��f��K^��e�f�g��{��R�*�/�2����+]��G�*��;X���o���sZ��2-X�����2�� �
/2�^�9t��2��*k�i�'�^��v�������	Z��,�e�=�ݭª E��:3�[������Ԙ�os�K]��5��Lg;���Sr��p+����tq}��Cթs�q�6B*I�`T�f�O]i).�3�|y�zU�Ǟ��V�%�N��}�Q�xb\?�C׬��YRL�O� ��M�+��@�o���z���SMx�h�i��L�	Fa�	*Vizqt�ňi?��/�.+Ce�1�������H�'�?\^�m�S�2Z`���qG�k1qDH0�j	 
t���Ul����x�G�%ޚ����D'j�)?���c���t�y��7@����g�3�;r�%|<��݉ ��F�|`�+��	��H��ط��X�_�ejB���B�\:V�W?�t�jV�=�2s{{ ���H��޻dG�2�Ӛ�!��W]��K�rPo*31��b5�!ŀ����5^��<^!���ӽ6}�k�w6�~+��.˟܊f>C�>��J�-j@0~C�"O��"P1�%�^26��{g5򞌃�$O{�{�뷯�/`��Yi$��	�6�m|)H��x�H�|x�YH��Ԓì��8WY��լy�F��'��F��-��h<~�����w��E��?�j�c^
\��D����>�<0��W0�m���o��~��y�]'�$�]����*ӳ&ۀ�q}�c�C,�R� ,�x&��x�k�8��9�3��J��V�˺�A���4�wFTDZ�+���h���g����Ǝ0���Z���KhS	��|:��I\��@���c2Ȗ5�L!4՞쿿lca��dϪ�D_0N���A~�s�����,����Ǥ�����������2a��i��C��4�@/`�Bj��<m��
|�^v\�!�㷴T/�1�O�Iq��'-�{��u��ԕ}8Xv� 9^�	9s%�e:�d�>JDý�
���k�▷>���1N׭��&��#F{�׃U�%oP�>0ޱ���-x
����{Q@Y��<T9E�3g�6���Y�ޯ��x��h��>�G�x��qI��s]��M|�2�B��|�2�D�h�y0�)��������q@����u��YGR�q�U�n���@pE�g�y�աfP�sL�M�\N�C�ЭX���%�=��$9 Cc]��#��T2��P����֍�g	{�8�~�)_�s1�E�`ߘ]@n.O|��q���tf�ԆY�����C�R~�r&���	�s4�V���f>w��6�	��&�Yo�����{�#��<�[UT����ת,�t��r+�	(g0ܦka�Y��gfY<'�,������9:�Q�" �M1cp��)��߹�儦7gl��-���BK�w7��5���jw�`������NE��V����F���f�� ڻ���iv�����&��S9^��Bj|�5��.�۪'�27��Bؘ)���G͔�tj�F�ݛ9f&�=~y]�"z�{�jP��r����KY�O�d7����m�N�?B���}# ����+.�~�Z�w^�+N���q�Y1E���d���#KI4C�֥�у;��%c���u�Ly� qTʋ���������^h���ʾl������|4	��Π�����n���G�J�Ϫ�����#ʚr�%{��k4b���u�����	�b�_�B�����_ZV���ë�4����d�|U�d��K��L::^�-���F�(q,�."���;����9�^��ms�,_eV���hkw�*h��ǮwL�]��d���1��?6WZ�nKuW?(�����n���f�1~ҠJB]�i!U�iHz�71vl��oq�-�N�DHu��EX��K:��_�鬗�pi@��cE�r]�oe���cSǭ7,���2i��KyXD�.����F�؅=�{��y�c��B���j��Zv��Y.b� �9
��� #��^0q�4�N���u�j�P"��DZnzh҂:�|}M����xv࿷�_mh(Bj��y���M76��|�rщi�i�"rew�G��x���Ǧr�Ǫ��>x^�m�˞��iI� ��̦zL��_�{����~�{\~� ���]QN\�[�ͭѯ�N��Gq��{Iy��� �!��h�9�"�H�mϝ!X���-E�U���^��`;k@��F=�A�!ˀ����ҷ��p7,j5�Lg�jIH�|���S��YQuGYG�������^�{A��O���*�>F��h�CנcA��uG �A7@{\����oH������z���8��<:��Ī_����:]:1���apmd�|�^�Nf:�d�#{X ((����������U��0�7wds3���?%Q1	N/�K�G߅�>�2˭S�G7����X�U��Z�5�?��S%+_.����sH�&?��|�9+p���h�i���a��	�Ǯ�:`�
o{��z�H�[�C%Ț� xfV>����4�����
��%�����P�u����rvA� ��Q����.�;�4b1��D�ژ�l)�������	�.�5ܐkU�s�flX�PxjA�yڈ"�Q��R������$�ھZ�Ǭ�l��=�;8���r��
���:Hh�a�ԓ�$R���D!���� 
�"�c��?�ڀ�G��NU���G����Q��B�s&���3%�2���z���,Vz{}9�bm<�V�z���ݔ5�}ܨM��1!ZV	�:�~,!Յ��z�n��b"b�,��sI4b���4w��>��*[ ��������y�J���d����r���f !�����r�Ŵ�{�������g�P��]/Y�������z�2�nd$�"�=>���@�(�p{�+҅.u=O���7^������E�<#��:i����1�������BJY$0�ҵ'�ѯ(� )Cp�G����l�D�Z
���ڰ������Z^��=o�]�y��^�k~�E/�cS�����j1���L�H����"9w��>3��|q�Ō+>�[��a����Ȁ,�L46a����(��\���2���vJ���*J�ݨ����4�X}p�o=��Ǯ<3��g]1t��nz�8��G��Y�Wb4:���� 0��Q�[J��U�ø(m	IOmؾ)%��v�W �d7��J�����+�Ċ&���UX����Ύv��An��R&}�@Y�/R�O�7��Ś��إl��>�|�ȇx����TмP�9�@������u�~�z 9*�"�P���>A`�LRM��r̾qdJ]�N-�ٰ�euȅ��F:?�@o��#�Ͷw�ٗ�eg'Ɛ�w�K�?��(��K/���Ûk`z�O��B�6��'I���^�#TzkI��;��{�>Sԓ~'���ҧ�.zm�5;i���4�Y��dE|{l��@�Ů��� ���(��]�n�MB$qf(��%$t��&y�R���#�����:--�X��rZX�Z�N{.�>%� �G�)^�c�/X�2C�h��杻ޜ\?kb�w�� �"U7���$5U0��M�W<�p����b�o/�]f-�%xxtU������
 �Iq�Ģhg���D{ŭ��HA\�`�e^��ӠS � [D�LS����7����*'��F�z������;A������u��q�Q�M��[�D�d�jʷ&�+���NJ��yn؛��|���mK�U�t��d��:T��g8��Etz�<�<!�5��+Z�W蓢��=娎4ڧ����Xuzc��4�)ngvm�k����n,�ϘU.f>�i�>��TsVR�("�~�Q*�8-�@w� �x�I��Ĭ�>�q&����.���0e�P��.�R�|�%5�j�p��i�M�~���y��<b�av$X��������]�J��AE w�1��m�!���'��.Ĺ���Ό�ޤQ#����Xn��\rA�n�*��A/�������9�F�W(d��{���d��'��R�����L�@�V�p;��#)ҧ�I�5��%� ����ݍ9��Y��D���a뭖�PF�0��ˮ� �$��e�Xh�/���%�����D����gUpX��1��:�<'2E��҄�����o�)ҋl`��5� �����$�gmw<�&C��8j�����)1E�C�p]�-������Y�	���JAEU������
�I)LOY�@\x���<�xK�d�uM�d�@�Q. h����n
���*n9�Y���R~>9��eq+)p����?H��A�?�!���|+"Ej�s2P�A��i��?f�gF~�
�Pe%x*<�g�N��I`�F,�T� z{�vin�x�E������JI'��=s`@l'�`jTz�0��8�r�[��0�BƁ_�R���Ǌz�V|%-h��8��|�wV	=)���!O�YJ|',x����t�Z/�{��GQCl��p�E��sa6��,+���kKv ����G�!��T�@�;�Ys�n4�vށ�KER����9��%]��s:�ν���6V�j�f�*���*o�X�j�ٶ��b�����o-=�O}%"�xN�eOQw��	1��M�>s�EϹf�ぴݓATq0�-p���.����E�L�w����\z�A��ѯ"��v>�V]7�)�Ed�"_��$�{�Q�sq%1N���;ڇ�­Kb	�'�������s����/��ڳqpم�w�"����OK��&7���(�h�H���>��XK�ֲ��L�K�
�8�O7�k�R�,p��a5��$��V,|B�9BE��W���xc�߯�t����l~Мp=R8ٝ��ι�N�^~�{r~��<He���){�`���y�G�D��r�}"����A0��m ����!kG�����'�RPX���Q���#: ɵm�tmAA��_�u��!��jo� �#&�
���CqKK��P��c`d^8D�%����:�x�y��&f��_?�h*W�m�WY̢��O
*�M�."6��$u#{��\߳�i�GMO�\N�V�P!�p"���R��=��M,�v���F�S����`�'*��1d8߈��K��j�mR�ǎ�SY7w�!⬵WZ�O4m�`�;���k���(�Q�Z���MZu~yÐ >���#�~FM��4��Vg��:[��Z��넔��o%��� ������.���[ʇ�n����#j#�NKj'W�i�?���"��"�{�r��}� ��n2UN��|.�ǏF"s�pC��x��m�/z즳��{��B�CP�-� <O�*����M�>�,������|���.��d{�� ������  %na7[e6�Ѡ�P�����{��Zk�H�WCy_�������a�%�Ά�!AX^�l]��`�'ۥ����݂������ѱ�7��@J�E�Y�Yt!��\k`�ؼ�wt�u��7��ۃ�FVbGqt��N�&�WH�Z��P�f�Om����l�W��]\>�G�;=�	�kW��To(Z���>5���ݝ0���瑖��V����U�ĸ��K�BܺL����|���i�#
\�=�-�J�p𼮶��	Z�K���>|��V�1���V�V��#+>�p����e���T�@������|��(�K{٭?��t�9^�����H��T�uX#c�	F�a���3�r㪧"3�T_���e�LX]卵<9���E�
�b�,�&�h,�`M�Qt�ɵ�Yr͉%WͶ�c:�F���[X���Q(���@���d����T�����=6_d���׏��"��^�\ �D!`��5�-l���Ȕ�,�j��-��� �+"A	+��,GYM�����؞T���5�υO���rL��@"0�C *˿�� ��B��L�^��V����c��7�4�"��x���ĸ�B=���^�D�1�Z}Kr^�4�i�^S}m�L��0��%*ؗ�a�{Wz�l����!+6��̀f�.Z؟��)-��F?,�8�+`:8(;�l�vVv�����i�]l a<�h�O[��Dk g�Xag�#%ee�呃���]O�{!@�8�Y��v���u�x�g���t�r�c�Sz��8�z/�Ki蔹C[���h���������&{C5x�r�t�2�#;�C�+S���R�y� ��pX?�F�����)�ш���$���T�vƃ�8X�)i����/ P�[��P�o3���ӥi��$^�t;����K��T�,��\)��|r����PX�9ڑ�a)ՒdM�yL�[��yzA������v���<_��)��I�2f$�}����'���*$kh9؉�L6uö��j/^�z���:��`E ��nxR��_���X�b�	��PRDع;��2{���u|�d�R��+�cBk����,���ێ�y"�������,�w��+���ӱ
%�#k�q1y��}���$��"��vڎ�!y�r/!?�p<L<S�g����|5��|l����s �{��`
.,�^�F�cx@͏׈�<� W���*i/ed�ſE��ސz5�p���4��d�c�{�#��G�[�愲8��f���i5-� PC�S�:���7E�Φ�O<��7A�>�#��/��DN3�;�:K��m�+c[
�l*Ju�oIB%3���WLN���WB�;o�%y��|�4�ar��}�������-��w(=���<摠'�"�]QiSv��1H8�c��h�>cQ�,��`�&A���^�K"�pK]��n�4j�����4+۝��B��8[���V�����`�d�=PY�������If�d �ξm����_0�P������#�N��H��E
XNAs��}��y����4���"�Y$�T�Tb1��խbJɴ� �W�S�󈦍�u������ؔڋ)T�����,ζ ��}{DxX�0�Q�h��B���e��֜P27���G9�v֪��hn����FH��B��_��nڿ^M�=���]q�3i����5�4�r)�b��G��-��x��0���^A\�����5~��[��ӯ�.7+��h{�|�O�qw��3r�D����qo�zn�9�q�0��O����w����*�i�f��k��a��p
�L������nt��=��}����Thϊ^�+-��Ӭ&�im��79��v�;D0RS������ս˾I�])�﷚�����08�����8��q��x��:PSŁ�@|�M!��We�|���N��[i�����Szp���&_��l��*�c�(��{����߭��oE��x��b��E۽=���E!��U��ºC�]0w�����a���v��84��ˏ�X�ҒR���\��;��Xtpt��LF�ܿ7,�����D�5Y�(�	!�����c�lH�X���@'|�:SS���A���??<��p�T�� G��ek��`m!Z@����9$TȰ!XZ�}/���%�SA����of��>�3h?���Q
�4
��DH�]ǳ��3�zG>�ӟ`�[�'t���4	bW�;��+�,Qb�_�?�w��59���2&`�&xԄ�Ăz�#��o�C�4G�q.6~���ݑ�P���^/��J��VpL����d�����_]�$�شN�wUUa�oH�aMσ�c�@��r�r�c��W�������x��D��a/�ը�j�Q�>�R�ǣS�`�꾷a�E:��1n6�[�,����Y佝/0��Jy53�cyW�?��V� �2��a5��c�?�~�j�O
���fD�\.'] m�5���kI�aT�G�o~S�Y�4��4�'	ɂ�7�g]2j[�+p_��$�#�T���B��*���,=��R�#��C�U�;��@�@�F�ѕ�&'�������;���7 �1;�N��)��פ���u�
�<	����#�+��Jmx��/��
��s��Ƣ/�=���Uͻ���/v� o��X�����ݤ^������1Kr�j�؃�����6)+ ��f����hZ��c�V�c���������I��Ͼ���T�!A0�\M�Y5���9u�16G?���_mK��K�j0��|��k��v]�+V�)Fl�BV��`Pe���P
��9��W%��3{��d���Z	�t/�2�w�#ބ��ȅϻ�!����L{7��S	�H:vE!␟8P���E#���	�]	�i,� \@`6rU����\��g��񥛍$"�j�Ȧ��E�ڧR�&���_�e���NTU8��B�/˓M'U	�ɄU��t>F�=��h�B�����{	���%Z��eP:�l3�,���X�����ڟ�f��0t3Yp�X���/�1J�Ah�9B& ��a5#ķҞ�̤��W���{��l�%�B��}	�t�t�9=ޛY�!�muk.Qe� B�DR�8'>�t������l��k�1~{�+p��J�{���Q�U��v��]rT�`q�u�ŀv,^_��,H��b��).�䵡;��E!�ȣL����8���[���m݇�F0��GJC1!��?Ul�k�� �m��
��yӋ�OzcC��ն9�SHz�q���&���HL���U��}���) Q�y����q�%�Ģl\��n�៖s��0��K��/��-�M���Lj�"x��TR�w�xA��[IDg��D���6>�w�G�OV��n�>fW�L'��R"t���$�vN��7���U����~�B�a��%4�U\>�����ߞ�܏z�*��k�A4j.���cX�bF�N4��4eꑑ��=�'	= �����5r�H)�l���K�{5ZC��iFbI���G�)P(O7�0���9�� R���#4'�V�?x�Yo��C�%�S��4+�gєs\k�?��3�R�f���8��Dy��L��ƺy&dU���Hço[�SR5� +����X���a0�L_���g�H�|����Z#;�F!; D���xY[aVO�k:
����=0W�3>zK��/�U�����G��N͆\+�Uµ|*i��e[c;zD��#�OIA��L��Q2�b"�y�_��f�Q�v������@[��u�ߺD`$|����,p������1%P���F�￞K
ď�j���X�����k�Wn�;}�2?���Wn[d�>8�~�s��=\̱�Y���e �1�A�3�䜷�D�W\&��^Ye��		t�p(j�Q����7�&md�7y�Et�$�w�"ˑp���e�n�mDF�~ϝ2Ē�2O�����r��\�;��?+�X�5bی�i(��.�3)�HGR�:���v1I�eNh�jm25�a�a�j䴿�h�%N�M'R�	OS�ճs=�(a�:�loޯփ�����"�� ^�T��=��&��d%TC��0 �%��b;����Ud	 Vݖ��/�Ԝ�JH���=�]�ߧ�w�y�z����N��1ƻC�>̒����/ ]^�;.��I҆ϴ/�ȸ��O^�Wׄn��F����M�Mb���ق7��Q?�U��b	�^�W'c7��8�KuoM^�5ZvH���LW_�Z;6�� ���x�;��*�?�D�:�W��9��f�s���.�͠V'յI�y��	%�K����o$~c�E�j�
{��[_�K� �f�h�xWb]5�٢D�"_�/����顟�Q�<�*IY�,׫H�
�ҝ���\1$H�Z5T�Շũ���!�z[=��Ų4����0YH;�f��$���8���B_OY27�S��IS� ��b^�}?�щ�#���֖����t���њ�Ѫ�`+���eI�/I�s@Vo��З����i�G�IgN_�����d�!)v	Z����jZ�֭,��^ܭw�)@��4����h-�2�����Q_�3�]���d�n�v�/�KU���I23]��K�a����<|�>�d	��t�`��2x�#
���t�W;X��H�5���$d6��w��������c��3�6��Xx+Ts���48wb w��,�*����%�M���^]�6��T(�˴#��V�o�mt_���z���SkQT���I��D�@�ӂ"�z��J��nOR���K'?���6>C$U�ڎ�$���9�G�/���D?�WɻW8Y&�^��=K���g<��B�jQ��C@��rUD���l���?�p�Î%���x�BгJ9%��L#.���{g�\����\��v���:���������$��|���gg-l�����v�W��h��G=�S�:���e��	��ҸyHY�2�9��t@��:�I�l0�9G����71H�i�����9����O����z�*w
���i/:o�����9�e�YNaӉ���Bzʼ�7�����uA/��|98|���>H������W$�j�K��W���R�	h@�������L�;�Ni������ �@2s9|i6�99\����)��n��0a([�Ɵ���C�~���B?�(�!��F̙@G�G��u�)�*�͈~R�����=�8�,b}���|"c^)S��g���^
�h W�4A ��dN��kr�,���&���$j��dF!�Q��E�*_c�٘ZS�c�E�$R���[.�K:<����P&��7Z���ß�'�#�e[�2�|e�>��m���(�Hr=BK��5�NZ]�F��|�f�g -α�Si�i���:r�<MXə^,��j�yNC�����lClg�j$��rC�$�r`�,V->0��F^��f�u-��e�0�2�_�3_6\H#�%'K)��R`*>�YmgY�2ܞY���7�.th�ik��\H��P6\+68��:�[�<��]�
��P0� �����$��f����N�U��G0� �����;1AW�pY]V`���`qg������@��vy�����+��̓�����>�E����Jg\���WS�f�&mL��~'�2f�q7�����.	O��y��Z����it۞'m�#ɣ���{l�A�	�N�����s'yPz3��x�����k��A�|��3R��ȣwʋ�� �[�����SE>.c�Q��v.筡��C��V�|��=�=E�\(X!Ux��o��`I��@*4��y��L�ă	^"��}��!�;�aVC�A)\�ۆ����d�4}�YS~Ρ�Ȕ�zR�6<j*�M2�3�[��5<Mb����ν�O�]��b6+��ve+�`x�bM����l�C�c��܃����}v�S�����L�=Q�Ge���7�R0���Mο����m�k2<��\#�(��ZL�LT������<E��O���F�_j�a��aC}���9�Ks�p�4Hc��^�-�������Ƴ�⑐n
]��$Ч)'��@<���yP5�FN8���{�ٴm��k��>��W��k�/��> 4}�җl~�� |Ͳ3Z[�P���K����*�p#`����Ɔ�b����2m��aӟ�ms��B���^[���}��c �h��|���kq<g�	��w�5H썿��CՃE/~�<��iҿ�EK�$�5���V�0�A"���'�%�Rd���ՎZ�S�V^~AM�ICL�5�e�U-�p�-�W��=�Oy�R+��������a����MQ��A��s�j>2�a�q�\�T���_���wzYr��n���54�DF�*���"�q�ؾ�`G��e/"1[y��>N�I1g�BaK�p�6R����uOrp���V��O����Ts�?��X}=4rqYK�%�<�c��΋] 2m/��������Ndl�ri@��P���\ �(�w��p�4�m ��Hyw0�����D��*qeeG���5s?��W���ɖ���Z�ü��ڋ?�J~���.5�Ap�&��6��'�+]��'݃r�.Il��s����B�t*���b�/����xomE��Ee��Zu���G�R��ƅ�rFgg �XX���5qf��yE��!��Z���F�w�L����]F,}���|㊕�mG���r����?=r�V4'��y}��:�5���=�.+Ӕb�)ـ驸�ΜNHzq� �E�j�A8/yf��=5����%����u�[%/�v[!�h��̐���Ե��H?��m"b����ka�u�Y�er<NZ����KV����󫋳r��fq��
�m�:��-�P��	��× �X�wKðoD��0@�U��q�.~j��Jt1�܉l��t��-v�<����x��.��'���uxN2h�\���fY'�=E�[�g�n{qj��y��q�M�|B��\��r������_��0%�B���T����ۇA��C*7Q�7�;m���c���('�()7~V~�?���.n`���b������͡�������*�f�45�Z8}�O���0��d
٭#��DՖ�	�*(jI��i�ԇ�`�sc��7N�H�X?q�����m�)���z�˴W�zx�\�-�2Y[R�?��sl��6�fA�1�j~�=ƍ�[��kZ�����9
�z*Ї.3��F�J�M^����'lb�~y�4���fc����5a!t��eQ�KS?�5�"�Vr��r�iv�3�'K��=Į G�8��+clTԧ�r}4��hz�f�Q�nVf<�rn��n2V?�S�%�}Њ�s�{���\+�TqV���`�-���e:=8�7�qfKD;g\�	�ɜ߉�s�0�[/��c�߸%"�m*rH�a\	OOn��K�[ H�[fu�������?�+Cx�no�̺�
�`�s������x۠�Ńi�b�=7�k����� ?��7�����ɞ��B�;�@QP#�$4�;Yo׵��ͳw7q8Uq_�w�SW����`r��,���ޱ��/LF���*���N���.a#Bb:�/ã�Ե���F �c1�&7<���gJD� �	���P6�7O��J�r�vͤ��豩�X$�GA*��F���.7���S��G�l�l�B�$��T��Ö[��1$�1	�y�e��t���H��1 ����Pp�'؎S�d� ��O��::��Q(:7�9�P0�.ߌ�M齏Jh��_������^�kgҒ4[�,����?qOv�t���"� �f��64|w�[m2�N�!�Ǧ.�aiI��RE��&3h)-�ZR��F|�*���ϹX�a$< be��v�T|͓"[�+���x���-5�%�d4�m8��������#�o�{���)[�Ւ��+�~Ux~�̀=UtXZ�OxN&X��6ks�П��K9���1u�����Z&��s�����pFm� 0k������.����xB5@q����F] �໷�%�Y�E#'K ��.r_��[��Q��3{}'�!�w�wR�"�Q���^?F@����ӹ�-�쓌h)R(Y
Q[ڕT�Hb���L�y���A�iz�7���I�YbR2p�c���L٠t��0
�����9SRppX�J5`HO�V*DĠ�Gi�l
�D^Y&Q���v}k�N�'�D��#�������o�s�XvB�h}�>�D�/�S���d��qz����X��i�l'̧JR��ʲ���e��?��t0�K���繱�v��A��N�41�6��<�>���
u�!o��:�^��ՍlDʢvG=�!N�Z���9cQ)���kӝ��+𵍠,C�(0{�Pj�� sH��73�~�_�ެ�y�9�ǫ�,�a�&�}��N{~��b���V`V�ٛ�7����;��4��b4��˶�V���+�ix�ܓ��Ǥ�����F�lł�阖	:���$"p�s]/�ȐoU���V�t� �Z�ě�k�&gF ��sv]0�K�l!�~,����ؼ�XO�,���:鎚�'ъ�s�'�0�&5M+�ײ���]c��yPߐ����vV߇5��j�E\<6u�C-�Qdv�_J;-38uB�I����?o4ۍ�(�x@��)M�w�h�P����#W	܌���g��r������ӎ�4�C����ه�1��vK~�iR��?TiY�fl�sg�=�SK(�]���'G�h�oH��>�Ǘ:(�!�R�I���@SwC����i5Њ{�,�ݛ}3�,m��'F��Ţ��I7�7�h�"F%��%�d��~I��^�O��{P��I=�5��yH*�b�!)	^m�z��������i�O�=�k� ��z�X���$�6욣Ì7�%�#�CO��`�V�X�T3�۹c�p���t�-9st[��~O���j9E��۪m�f+�=�)VJT8������
�r���Ȑ��d\�V�G�!�\G?���L2P�~��vB'�7m�S�["9��9OU�
�K�vUѸ�g��H���~ϔ�+J�͚��ȡj��O����C��dfL3�5b/�T�5Q{�Eh�)�f��@�i}�^�$��co� �����zR˰�®ӌ���;��e�1&p�k��2j�q��;�x��|ar��X����{�cԽ��b�ـ)�R��fL���nw����ꀷ�|�F+$ײ�Z��B�/y�<L%�%x���V�ȆS��,M���[��m����C��^cD�BA"#�K�p P���3g���T�	��{p��	�����7��2g?���^�����d���7�τ�=����&�ń� �����h��+A8�S���r*^b�K|����)��ȯ���{I���f304�o�;��������}�؄<?�� ����ğ��1�,�|��Zn�XzpL �@�#����+�4��j�-ىE����o����.�����unOP�������6Ԋ�D2��1	�w�X����:�Z�=�s�!�`��%���}�#�Za5eD�u#��6�+db��1�KsV�I����#D�D!��,=���z+��V��O=v6�9&�{ ՗D�`���XE��.y����_*uå�,m���		z��{l�_�l+[��XW4�d%�d�{7��=)e +�VP:t&�[����3P�Q+ӒȊ}����\�%et^�����A���ſ�OJ�K�W��)�>�|4�.����P�SW̪/ė��ɵP?X�HW�_�-��3��$q8�r�r߈��aF��!�ɿ6�sϘX���g�A1�x�yc�nn(<A����^��O]bl�⚧:���Ǹ^xC���1̌��MǤ�/_z�꩏�X`y������ңw�}KTD�~X�b�J���Ol�����pQ�&��8�Rd�&�	�y����ך~��'����Iz\ͭ� �ླ�Ե!�����h�^��4��u� ���]Ő�K��;�-L�gX��yr�3-���J�uY�Jɡ1,1�g�5�ė,�I��jmz���7~�rdL��Csx����4�D�u���v���,aK�ǁ�t�z{�D*KK� �B9ۚ����A�������LX0g�.��*�K��5�8���u���ˎ�ڒT��p��C�8��.�O�2�;=��X�H��������(���t�c*e��G���|w����//-<CV��ϙjg��Иo�f���/���:O g�m��k߬zX��,ϣ�0�ES
0TH�A��ر0�hvX�E�uٚ򛬫��ܽ�`>]`� 
�4��J�]Ⱥ6�	�,�W!
�6�%)������\G�x�N�Ў��N]֓�c�%A{b�%xa�7��V�oV����JJNv|pN�$�X?`�5�k����{)�B��fjY�>7����J|�D���f0�%�H��C0(]�?,���N���I9kG�٧�M���~�SS�@٬?4^��迒cR�E��ƶ��ȳ���ߠd���'���>��_��,HE����9r㾆o���i���]��#^R�R��E���#�LEm Z���K�*��V�	�9����F�#3�P��9�
:�(�����u;��9]j���\S=;o�0�������Ҳ����V��s,�(��<�~�nپ��$#h���꥘o�jW`��$���5��=p��-���2��?Pd�z^�����0�/��["[��2��7���/r��ƹnQ�k%�`���� ��7�{5U���C����m���.�e.����K��F�rc�x������(�l��P��p�|�&3�C��� �&ZQl�Ȩ9���~x7�W��М�4���+B`$4j��c�ut=	'�@4�C�}�m��cWw����PI�J0(}(�!�-�{F'4i���_�6�����7;(��4����F�>&�8�D4<.�lO3��߰Z�뻀��Г�^�sTr�B��L���b���V���!`�<��Է�g���g��c{��o5�0���cqn��<��KT�}X!��ۏ
cX�t�A1�=1w�_����A�s@��LTc�`��0
�ԫQ���}�l���{�j�M5��m����Y�K|�K)<$������t�_�޴�dK�s,�
-���^KA�mi���ܕ�T�9���?	[P>A�az��y���L��8��~��J�� 4C�];7��#���oF�C�0{�<���ɬ���b���T�U��yӑ���μ��+�pI�p��ʫxe�Ny�o4�� ��CO�F�h��4����$FW[�!G�Uۙ�E���e���yޥ��|�Ƌ��h[���O���C���׾$C#^�l�4�A=���:�w�O�ɦ�ޭ���6d�] �2��Y�YYnW�(}N��+.��m����}�v6�Ji��՜'���p�q�@�{�a�I�����E(G�/�Ǧ�:�eŕT0�m�Q�o3���^�/��o��I�"�~�:��L�Z?�TNT\�k~��<0rLv�nR��^̫��3[�o|����д��S�r\/.�jϮ?�"2�l	q��R����6L2kS������^�5�� �"�P ����|�zX�� ��d�U4a["�2T�"�� W�fβ3���8��+)��&H�,����(��щl\����̦���%��y$�c�j-��xP�.}(�<ֳ�왷퍃��R�ع�I��bM�j��_A�6�����
��g� ���G���J�P��0eO�ݰ�o�B���u렕.K�����?�95f3��$B����	'�Dv��