// soc_system.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,       //      alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,      //                                 .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,     //                                 .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid, //                                 .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,    //                                 .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,    //                                 .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,         //                                 .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,         //                                 .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,         //                                 .vid_v
		input  wire        clk_clk,                                   //                              clk.clk
		output wire        clk_sdram_clk,                             //                        clk_sdram.clk
		output wire        clk_vga_clk,                               //                          clk_vga.clk
		output wire        d8m_xclkin_clk,                            //                       d8m_xclkin.clk
		output wire        hps_0_h2f_reset_reset_n,                   //                  hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK,     //                     hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,       //                                 .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,       //                                 .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,       //                                 .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,       //                                 .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,       //                                 .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,       //                                 .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,        //                                 .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL,     //                                 .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL,     //                                 .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK,     //                                 .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,       //                                 .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,       //                                 .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,       //                                 .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,         //                                 .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,         //                                 .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,         //                                 .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,         //                                 .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,         //                                 .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,         //                                 .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,         //                                 .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,          //                                 .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,          //                                 .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,         //                                 .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,          //                                 .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,          //                                 .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,          //                                 .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,          //                                 .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,          //                                 .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,          //                                 .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,          //                                 .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,          //                                 .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,          //                                 .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,          //                                 .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,         //                                 .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,         //                                 .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,         //                                 .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,         //                                 .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,        //                                 .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,       //                                 .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,       //                                 .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,        //                                 .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,         //                                 .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,         //                                 .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,         //                                 .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,         //                                 .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,         //                                 .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,         //                                 .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,      //                                 .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,      //                                 .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,      //                                 .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,      //                                 .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,      //                                 .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,      //                                 .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,      //                                 .hps_io_gpio_inst_GPIO61
		inout  wire        i2c_opencores_camera_export_scl_pad_io,    //      i2c_opencores_camera_export.scl_pad_io
		inout  wire        i2c_opencores_camera_export_sda_pad_io,    //                                 .sda_pad_io
		inout  wire        i2c_opencores_mipi_export_scl_pad_io,      //        i2c_opencores_mipi_export.scl_pad_io
		inout  wire        i2c_opencores_mipi_export_sda_pad_io,      //                                 .sda_pad_io
		input  wire [3:0]  key_external_connection_export,            //          key_external_connection.export
		output wire [9:0]  led_external_connection_export,            //          led_external_connection.export
		output wire [14:0] memory_mem_a,                              //                           memory.mem_a
		output wire [2:0]  memory_mem_ba,                             //                                 .mem_ba
		output wire        memory_mem_ck,                             //                                 .mem_ck
		output wire        memory_mem_ck_n,                           //                                 .mem_ck_n
		output wire        memory_mem_cke,                            //                                 .mem_cke
		output wire        memory_mem_cs_n,                           //                                 .mem_cs_n
		output wire        memory_mem_ras_n,                          //                                 .mem_ras_n
		output wire        memory_mem_cas_n,                          //                                 .mem_cas_n
		output wire        memory_mem_we_n,                           //                                 .mem_we_n
		output wire        memory_mem_reset_n,                        //                                 .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                             //                                 .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                            //                                 .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                          //                                 .mem_dqs_n
		output wire        memory_mem_odt,                            //                                 .mem_odt
		output wire [3:0]  memory_mem_dm,                             //                                 .mem_dm
		input  wire        memory_oct_rzqin,                          //                                 .oct_rzqin
		output wire        mipi_pwdn_n_external_connection_export,    //  mipi_pwdn_n_external_connection.export
		output wire        mipi_reset_n_external_connection_export,   // mipi_reset_n_external_connection.export
		input  wire        reset_reset_n,                             //                            reset.reset_n
		output wire [12:0] sdram_wire_addr,                           //                       sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                             //                                 .ba
		output wire        sdram_wire_cas_n,                          //                                 .cas_n
		output wire        sdram_wire_cke,                            //                                 .cke
		output wire        sdram_wire_cs_n,                           //                                 .cs_n
		inout  wire [15:0] sdram_wire_dq,                             //                                 .dq
		output wire [1:0]  sdram_wire_dqm,                            //                                 .dqm
		output wire        sdram_wire_ras_n,                          //                                 .ras_n
		output wire        sdram_wire_we_n,                           //                                 .we_n
		input  wire [9:0]  sw_external_connection_export,             //           sw_external_connection.export
		input  wire [11:0] terasic_camera_0_conduit_end_D,            //     terasic_camera_0_conduit_end.D
		input  wire        terasic_camera_0_conduit_end_FVAL,         //                                 .FVAL
		input  wire        terasic_camera_0_conduit_end_LVAL,         //                                 .LVAL
		input  wire        terasic_camera_0_conduit_end_PIXCLK        //                                 .PIXCLK
	);

	wire          video_csc_0_avalon_csc_source_valid;                                          // video_csc_0:stream_out_valid -> video_dma_controller_0:stream_valid
	wire    [7:0] video_csc_0_avalon_csc_source_data;                                           // video_csc_0:stream_out_data -> video_dma_controller_0:stream_data
	wire          video_csc_0_avalon_csc_source_ready;                                          // video_dma_controller_0:stream_ready -> video_csc_0:stream_out_ready
	wire          video_csc_0_avalon_csc_source_startofpacket;                                  // video_csc_0:stream_out_startofpacket -> video_dma_controller_0:stream_startofpacket
	wire          video_csc_0_avalon_csc_source_endofpacket;                                    // video_csc_0:stream_out_endofpacket -> video_dma_controller_0:stream_endofpacket
	wire          terasic_camera_0_avalon_streaming_source_valid;                               // TERASIC_CAMERA_0:st_valid -> alt_vip_cl_clp_1:din_valid
	wire   [23:0] terasic_camera_0_avalon_streaming_source_data;                                // TERASIC_CAMERA_0:st_data -> alt_vip_cl_clp_1:din_data
	wire          terasic_camera_0_avalon_streaming_source_ready;                               // alt_vip_cl_clp_1:din_ready -> TERASIC_CAMERA_0:st_ready
	wire          terasic_camera_0_avalon_streaming_source_startofpacket;                       // TERASIC_CAMERA_0:st_sop -> alt_vip_cl_clp_1:din_startofpacket
	wire          terasic_camera_0_avalon_streaming_source_endofpacket;                         // TERASIC_CAMERA_0:st_eop -> alt_vip_cl_clp_1:din_endofpacket
	wire          alt_vip_vfr_vga_avalon_streaming_source_valid;                                // alt_vip_vfr_vga:dout_valid -> alt_vip_cpr_0:din0_valid
	wire   [31:0] alt_vip_vfr_vga_avalon_streaming_source_data;                                 // alt_vip_vfr_vga:dout_data -> alt_vip_cpr_0:din0_data
	wire          alt_vip_vfr_vga_avalon_streaming_source_ready;                                // alt_vip_cpr_0:din0_ready -> alt_vip_vfr_vga:dout_ready
	wire          alt_vip_vfr_vga_avalon_streaming_source_startofpacket;                        // alt_vip_vfr_vga:dout_startofpacket -> alt_vip_cpr_0:din0_startofpacket
	wire          alt_vip_vfr_vga_avalon_streaming_source_endofpacket;                          // alt_vip_vfr_vga:dout_endofpacket -> alt_vip_cpr_0:din0_endofpacket
	wire          alt_vip_cl_clp_1_dout_valid;                                                  // alt_vip_cl_clp_1:dout_valid -> alt_vip_cl_scl_0:din_valid
	wire   [23:0] alt_vip_cl_clp_1_dout_data;                                                   // alt_vip_cl_clp_1:dout_data -> alt_vip_cl_scl_0:din_data
	wire          alt_vip_cl_clp_1_dout_ready;                                                  // alt_vip_cl_scl_0:din_ready -> alt_vip_cl_clp_1:dout_ready
	wire          alt_vip_cl_clp_1_dout_startofpacket;                                          // alt_vip_cl_clp_1:dout_startofpacket -> alt_vip_cl_scl_0:din_startofpacket
	wire          alt_vip_cl_clp_1_dout_endofpacket;                                            // alt_vip_cl_clp_1:dout_endofpacket -> alt_vip_cl_scl_0:din_endofpacket
	wire          alt_vip_cl_scl_0_dout_valid;                                                  // alt_vip_cl_scl_0:dout_valid -> alt_vip_vfb_0:din_valid
	wire   [23:0] alt_vip_cl_scl_0_dout_data;                                                   // alt_vip_cl_scl_0:dout_data -> alt_vip_vfb_0:din_data
	wire          alt_vip_cl_scl_0_dout_ready;                                                  // alt_vip_vfb_0:din_ready -> alt_vip_cl_scl_0:dout_ready
	wire          alt_vip_cl_scl_0_dout_startofpacket;                                          // alt_vip_cl_scl_0:dout_startofpacket -> alt_vip_vfb_0:din_startofpacket
	wire          alt_vip_cl_scl_0_dout_endofpacket;                                            // alt_vip_cl_scl_0:dout_endofpacket -> alt_vip_vfb_0:din_endofpacket
	wire          alt_vip_mix_0_dout_valid;                                                     // alt_vip_mix_0:dout_valid -> alt_vip_itc_0:is_valid
	wire   [23:0] alt_vip_mix_0_dout_data;                                                      // alt_vip_mix_0:dout_data -> alt_vip_itc_0:is_data
	wire          alt_vip_mix_0_dout_ready;                                                     // alt_vip_itc_0:is_ready -> alt_vip_mix_0:dout_ready
	wire          alt_vip_mix_0_dout_startofpacket;                                             // alt_vip_mix_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire          alt_vip_mix_0_dout_endofpacket;                                               // alt_vip_mix_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire          alt_vip_vfb_0_dout_valid;                                                     // alt_vip_vfb_0:dout_valid -> alt_vip_cpr_2:din0_valid
	wire   [23:0] alt_vip_vfb_0_dout_data;                                                      // alt_vip_vfb_0:dout_data -> alt_vip_cpr_2:din0_data
	wire          alt_vip_vfb_0_dout_ready;                                                     // alt_vip_cpr_2:din0_ready -> alt_vip_vfb_0:dout_ready
	wire          alt_vip_vfb_0_dout_startofpacket;                                             // alt_vip_vfb_0:dout_startofpacket -> alt_vip_cpr_2:din0_startofpacket
	wire          alt_vip_vfb_0_dout_endofpacket;                                               // alt_vip_vfb_0:dout_endofpacket -> alt_vip_cpr_2:din0_endofpacket
	wire          alt_vip_cl_tpg_0_dout_valid;                                                  // alt_vip_cl_tpg_0:dout_valid -> alt_vip_mix_0:din_2_valid
	wire   [23:0] alt_vip_cl_tpg_0_dout_data;                                                   // alt_vip_cl_tpg_0:dout_data -> alt_vip_mix_0:din_2_data
	wire          alt_vip_cl_tpg_0_dout_ready;                                                  // alt_vip_mix_0:din_2_ready -> alt_vip_cl_tpg_0:dout_ready
	wire          alt_vip_cl_tpg_0_dout_startofpacket;                                          // alt_vip_cl_tpg_0:dout_startofpacket -> alt_vip_mix_0:din_2_startofpacket
	wire          alt_vip_cl_tpg_0_dout_endofpacket;                                            // alt_vip_cl_tpg_0:dout_endofpacket -> alt_vip_mix_0:din_2_endofpacket
	wire          alt_vip_cpr_2_dout0_valid;                                                    // alt_vip_cpr_2:dout0_valid -> alt_vip_cpr_1:din0_valid
	wire   [23:0] alt_vip_cpr_2_dout0_data;                                                     // alt_vip_cpr_2:dout0_data -> alt_vip_cpr_1:din0_data
	wire          alt_vip_cpr_2_dout0_ready;                                                    // alt_vip_cpr_1:din0_ready -> alt_vip_cpr_2:dout0_ready
	wire          alt_vip_cpr_2_dout0_startofpacket;                                            // alt_vip_cpr_2:dout0_startofpacket -> alt_vip_cpr_1:din0_startofpacket
	wire          alt_vip_cpr_2_dout0_endofpacket;                                              // alt_vip_cpr_2:dout0_endofpacket -> alt_vip_cpr_1:din0_endofpacket
	wire          alt_vip_cpr_0_dout0_valid;                                                    // alt_vip_cpr_0:dout0_valid -> alt_vip_mix_0:din_0_valid
	wire   [23:0] alt_vip_cpr_0_dout0_data;                                                     // alt_vip_cpr_0:dout0_data -> alt_vip_mix_0:din_0_data
	wire          alt_vip_cpr_0_dout0_ready;                                                    // alt_vip_mix_0:din_0_ready -> alt_vip_cpr_0:dout0_ready
	wire          alt_vip_cpr_0_dout0_startofpacket;                                            // alt_vip_cpr_0:dout0_startofpacket -> alt_vip_mix_0:din_0_startofpacket
	wire          alt_vip_cpr_0_dout0_endofpacket;                                              // alt_vip_cpr_0:dout0_endofpacket -> alt_vip_mix_0:din_0_endofpacket
	wire          alt_vip_cpr_1_dout0_valid;                                                    // alt_vip_cpr_1:dout0_valid -> alt_vip_mix_0:din_1_valid
	wire   [23:0] alt_vip_cpr_1_dout0_data;                                                     // alt_vip_cpr_1:dout0_data -> alt_vip_mix_0:din_1_data
	wire          alt_vip_cpr_1_dout0_ready;                                                    // alt_vip_mix_0:din_1_ready -> alt_vip_cpr_1:dout0_ready
	wire          alt_vip_cpr_1_dout0_startofpacket;                                            // alt_vip_cpr_1:dout0_startofpacket -> alt_vip_mix_0:din_1_startofpacket
	wire          alt_vip_cpr_1_dout0_endofpacket;                                              // alt_vip_cpr_1:dout0_endofpacket -> alt_vip_mix_0:din_1_endofpacket
	wire          alt_vip_cpr_2_dout1_valid;                                                    // alt_vip_cpr_2:dout1_valid -> st_adapter_0:in_0_valid
	wire   [23:0] alt_vip_cpr_2_dout1_data;                                                     // alt_vip_cpr_2:dout1_data -> st_adapter_0:in_0_data
	wire          alt_vip_cpr_2_dout1_ready;                                                    // st_adapter_0:in_0_ready -> alt_vip_cpr_2:dout1_ready
	wire          alt_vip_cpr_2_dout1_startofpacket;                                            // alt_vip_cpr_2:dout1_startofpacket -> st_adapter_0:in_0_startofpacket
	wire          alt_vip_cpr_2_dout1_endofpacket;                                              // alt_vip_cpr_2:dout1_endofpacket -> st_adapter_0:in_0_endofpacket
	wire          st_adapter_0_out_0_valid;                                                     // st_adapter_0:out_0_valid -> video_csc_0:stream_in_valid
	wire   [23:0] st_adapter_0_out_0_data;                                                      // st_adapter_0:out_0_data -> video_csc_0:stream_in_data
	wire          st_adapter_0_out_0_ready;                                                     // video_csc_0:stream_in_ready -> st_adapter_0:out_0_ready
	wire          st_adapter_0_out_0_startofpacket;                                             // st_adapter_0:out_0_startofpacket -> video_csc_0:stream_in_startofpacket
	wire          st_adapter_0_out_0_endofpacket;                                               // st_adapter_0:out_0_endofpacket -> video_csc_0:stream_in_endofpacket
	wire          pll_0_outclk0_clk;                                                            // pll_0:outclk_0 -> [TERASIC_CAMERA_0:clk, alt_vip_cl_clp_1:main_clock, alt_vip_cl_scl_0:main_clock, alt_vip_cl_tpg_0:main_clock, alt_vip_cpr_0:clock, alt_vip_cpr_1:clock, alt_vip_cpr_2:clock, alt_vip_itc_0:is_clk, alt_vip_mix_0:clock, alt_vip_vfb_0:clock, alt_vip_vfr_vga:clock, alt_vip_vfr_vga:master_clock, mm_interconnect_0:pll_0_outclk0_clk, mm_interconnect_1:pll_0_outclk0_clk, mm_interconnect_2:pll_0_outclk0_clk, mm_interconnect_3:pll_0_outclk0_clk, onchip_memory:clk, rst_controller:clk, sdram:clk, st_adapter_0:in_clk_0_clk, video_csc_0:clk, video_dma_controller_0:clk]
	wire          video_dma_controller_0_avalon_dma_master_waitrequest;                         // mm_interconnect_0:video_dma_controller_0_avalon_dma_master_waitrequest -> video_dma_controller_0:master_waitrequest
	wire   [31:0] video_dma_controller_0_avalon_dma_master_address;                             // video_dma_controller_0:master_address -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_address
	wire          video_dma_controller_0_avalon_dma_master_write;                               // video_dma_controller_0:master_write -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_write
	wire    [7:0] video_dma_controller_0_avalon_dma_master_writedata;                           // video_dma_controller_0:master_writedata -> mm_interconnect_0:video_dma_controller_0_avalon_dma_master_writedata
	wire          mm_interconnect_0_onchip_memory_s1_chipselect;                                // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire   [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                                  // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire   [15:0] mm_interconnect_0_onchip_memory_s1_address;                                   // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire    [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                                // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire          mm_interconnect_0_onchip_memory_s1_write;                                     // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire   [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                                 // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire          mm_interconnect_0_onchip_memory_s1_clken;                                     // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire  [127:0] alt_vip_vfr_vga_avalon_master_readdata;                                       // mm_interconnect_1:alt_vip_vfr_vga_avalon_master_readdata -> alt_vip_vfr_vga:master_readdata
	wire          alt_vip_vfr_vga_avalon_master_waitrequest;                                    // mm_interconnect_1:alt_vip_vfr_vga_avalon_master_waitrequest -> alt_vip_vfr_vga:master_waitrequest
	wire   [31:0] alt_vip_vfr_vga_avalon_master_address;                                        // alt_vip_vfr_vga:master_address -> mm_interconnect_1:alt_vip_vfr_vga_avalon_master_address
	wire          alt_vip_vfr_vga_avalon_master_read;                                           // alt_vip_vfr_vga:master_read -> mm_interconnect_1:alt_vip_vfr_vga_avalon_master_read
	wire          alt_vip_vfr_vga_avalon_master_readdatavalid;                                  // mm_interconnect_1:alt_vip_vfr_vga_avalon_master_readdatavalid -> alt_vip_vfr_vga:master_readdatavalid
	wire    [5:0] alt_vip_vfr_vga_avalon_master_burstcount;                                     // alt_vip_vfr_vga:master_burstcount -> mm_interconnect_1:alt_vip_vfr_vga_avalon_master_burstcount
	wire   [31:0] master_secure_master_readdata;                                                // mm_interconnect_1:master_secure_master_readdata -> master_secure:master_readdata
	wire          master_secure_master_waitrequest;                                             // mm_interconnect_1:master_secure_master_waitrequest -> master_secure:master_waitrequest
	wire   [31:0] master_secure_master_address;                                                 // master_secure:master_address -> mm_interconnect_1:master_secure_master_address
	wire          master_secure_master_read;                                                    // master_secure:master_read -> mm_interconnect_1:master_secure_master_read
	wire    [3:0] master_secure_master_byteenable;                                              // master_secure:master_byteenable -> mm_interconnect_1:master_secure_master_byteenable
	wire          master_secure_master_readdatavalid;                                           // mm_interconnect_1:master_secure_master_readdatavalid -> master_secure:master_readdatavalid
	wire          master_secure_master_write;                                                   // master_secure:master_write -> mm_interconnect_1:master_secure_master_write
	wire   [31:0] master_secure_master_writedata;                                               // master_secure:master_writedata -> mm_interconnect_1:master_secure_master_writedata
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_awburst;                                // mm_interconnect_1:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [4:0] mm_interconnect_1_hps_0_f2h_axi_slave_awuser;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_arlen;                                  // mm_interconnect_1:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire   [15:0] mm_interconnect_1_hps_0_f2h_axi_slave_wstrb;                                  // mm_interconnect_1:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_wready;                                 // hps_0:f2h_WREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_wready
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_rid;                                    // hps_0:f2h_RID -> mm_interconnect_1:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_rready;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_awlen;                                  // mm_interconnect_1:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_wid;                                    // mm_interconnect_1:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_arcache;                                // mm_interconnect_1:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_wvalid;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire   [31:0] mm_interconnect_1_hps_0_f2h_axi_slave_araddr;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_arprot;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_awprot;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire  [127:0] mm_interconnect_1_hps_0_f2h_axi_slave_wdata;                                  // mm_interconnect_1:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_arvalid;                                // mm_interconnect_1:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_awcache;                                // mm_interconnect_1:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_arid;                                   // mm_interconnect_1:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_arlock;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_awlock;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire   [31:0] mm_interconnect_1_hps_0_f2h_axi_slave_awaddr;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_bresp;                                  // hps_0:f2h_BRESP -> mm_interconnect_1:hps_0_f2h_axi_slave_bresp
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_arready;                                // hps_0:f2h_ARREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_arready
	wire  [127:0] mm_interconnect_1_hps_0_f2h_axi_slave_rdata;                                  // hps_0:f2h_RDATA -> mm_interconnect_1:hps_0_f2h_axi_slave_rdata
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_awready;                                // hps_0:f2h_AWREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_awready
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_arburst;                                // mm_interconnect_1:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_arsize;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_bready;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_rlast;                                  // hps_0:f2h_RLAST -> mm_interconnect_1:hps_0_f2h_axi_slave_rlast
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_wlast;                                  // mm_interconnect_1:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_rresp;                                  // hps_0:f2h_RRESP -> mm_interconnect_1:hps_0_f2h_axi_slave_rresp
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_awid;                                   // mm_interconnect_1:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_bid;                                    // hps_0:f2h_BID -> mm_interconnect_1:hps_0_f2h_axi_slave_bid
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_bvalid;                                 // hps_0:f2h_BVALID -> mm_interconnect_1:hps_0_f2h_axi_slave_bvalid
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_awsize;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_awvalid;                                // mm_interconnect_1:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [4:0] mm_interconnect_1_hps_0_f2h_axi_slave_aruser;                                 // mm_interconnect_1:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_rvalid;                                 // hps_0:f2h_RVALID -> mm_interconnect_1:hps_0_f2h_axi_slave_rvalid
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                                 // hps_0:h2f_AWBURST -> mm_interconnect_2:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                                   // hps_0:h2f_ARLEN -> mm_interconnect_2:hps_0_h2f_axi_master_arlen
	wire    [7:0] hps_0_h2f_axi_master_wstrb;                                                   // hps_0:h2f_WSTRB -> mm_interconnect_2:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                                  // mm_interconnect_2:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                                     // mm_interconnect_2:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                                  // hps_0:h2f_RREADY -> mm_interconnect_2:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                                   // hps_0:h2f_AWLEN -> mm_interconnect_2:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                                     // hps_0:h2f_WID -> mm_interconnect_2:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                                 // hps_0:h2f_ARCACHE -> mm_interconnect_2:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                                  // hps_0:h2f_WVALID -> mm_interconnect_2:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                                  // hps_0:h2f_ARADDR -> mm_interconnect_2:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                                  // hps_0:h2f_ARPROT -> mm_interconnect_2:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                                  // hps_0:h2f_AWPROT -> mm_interconnect_2:hps_0_h2f_axi_master_awprot
	wire   [63:0] hps_0_h2f_axi_master_wdata;                                                   // hps_0:h2f_WDATA -> mm_interconnect_2:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                                 // hps_0:h2f_ARVALID -> mm_interconnect_2:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                                 // hps_0:h2f_AWCACHE -> mm_interconnect_2:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                                    // hps_0:h2f_ARID -> mm_interconnect_2:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                                  // hps_0:h2f_ARLOCK -> mm_interconnect_2:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                                  // hps_0:h2f_AWLOCK -> mm_interconnect_2:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                                  // hps_0:h2f_AWADDR -> mm_interconnect_2:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                                   // mm_interconnect_2:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                                 // mm_interconnect_2:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire   [63:0] hps_0_h2f_axi_master_rdata;                                                   // mm_interconnect_2:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                                 // mm_interconnect_2:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                                 // hps_0:h2f_ARBURST -> mm_interconnect_2:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                                  // hps_0:h2f_ARSIZE -> mm_interconnect_2:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                                  // hps_0:h2f_BREADY -> mm_interconnect_2:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                                   // mm_interconnect_2:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                                   // hps_0:h2f_WLAST -> mm_interconnect_2:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                                   // mm_interconnect_2:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                                    // hps_0:h2f_AWID -> mm_interconnect_2:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                                     // mm_interconnect_2:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                                  // mm_interconnect_2:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                                  // hps_0:h2f_AWSIZE -> mm_interconnect_2:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                                 // hps_0:h2f_AWVALID -> mm_interconnect_2:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                                  // mm_interconnect_2:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire          alt_vip_vfb_0_read_master_waitrequest;                                        // mm_interconnect_2:alt_vip_vfb_0_read_master_waitrequest -> alt_vip_vfb_0:read_master_av_waitrequest
	wire   [31:0] alt_vip_vfb_0_read_master_readdata;                                           // mm_interconnect_2:alt_vip_vfb_0_read_master_readdata -> alt_vip_vfb_0:read_master_av_readdata
	wire   [31:0] alt_vip_vfb_0_read_master_address;                                            // alt_vip_vfb_0:read_master_av_address -> mm_interconnect_2:alt_vip_vfb_0_read_master_address
	wire          alt_vip_vfb_0_read_master_read;                                               // alt_vip_vfb_0:read_master_av_read -> mm_interconnect_2:alt_vip_vfb_0_read_master_read
	wire          alt_vip_vfb_0_read_master_readdatavalid;                                      // mm_interconnect_2:alt_vip_vfb_0_read_master_readdatavalid -> alt_vip_vfb_0:read_master_av_readdatavalid
	wire    [2:0] alt_vip_vfb_0_read_master_burstcount;                                         // alt_vip_vfb_0:read_master_av_burstcount -> mm_interconnect_2:alt_vip_vfb_0_read_master_burstcount
	wire          alt_vip_vfb_0_write_master_waitrequest;                                       // mm_interconnect_2:alt_vip_vfb_0_write_master_waitrequest -> alt_vip_vfb_0:write_master_av_waitrequest
	wire   [31:0] alt_vip_vfb_0_write_master_address;                                           // alt_vip_vfb_0:write_master_av_address -> mm_interconnect_2:alt_vip_vfb_0_write_master_address
	wire          alt_vip_vfb_0_write_master_write;                                             // alt_vip_vfb_0:write_master_av_write -> mm_interconnect_2:alt_vip_vfb_0_write_master_write
	wire   [31:0] alt_vip_vfb_0_write_master_writedata;                                         // alt_vip_vfb_0:write_master_av_writedata -> mm_interconnect_2:alt_vip_vfb_0_write_master_writedata
	wire    [2:0] alt_vip_vfb_0_write_master_burstcount;                                        // alt_vip_vfb_0:write_master_av_burstcount -> mm_interconnect_2:alt_vip_vfb_0_write_master_burstcount
	wire          mm_interconnect_2_sdram_s1_chipselect;                                        // mm_interconnect_2:sdram_s1_chipselect -> sdram:az_cs
	wire   [15:0] mm_interconnect_2_sdram_s1_readdata;                                          // sdram:za_data -> mm_interconnect_2:sdram_s1_readdata
	wire          mm_interconnect_2_sdram_s1_waitrequest;                                       // sdram:za_waitrequest -> mm_interconnect_2:sdram_s1_waitrequest
	wire   [24:0] mm_interconnect_2_sdram_s1_address;                                           // mm_interconnect_2:sdram_s1_address -> sdram:az_addr
	wire          mm_interconnect_2_sdram_s1_read;                                              // mm_interconnect_2:sdram_s1_read -> sdram:az_rd_n
	wire    [1:0] mm_interconnect_2_sdram_s1_byteenable;                                        // mm_interconnect_2:sdram_s1_byteenable -> sdram:az_be_n
	wire          mm_interconnect_2_sdram_s1_readdatavalid;                                     // sdram:za_valid -> mm_interconnect_2:sdram_s1_readdatavalid
	wire          mm_interconnect_2_sdram_s1_write;                                             // mm_interconnect_2:sdram_s1_write -> sdram:az_wr_n
	wire   [15:0] mm_interconnect_2_sdram_s1_writedata;                                         // mm_interconnect_2:sdram_s1_writedata -> sdram:az_data
	wire          mm_interconnect_2_onchip_memory_s2_chipselect;                                // mm_interconnect_2:onchip_memory_s2_chipselect -> onchip_memory:chipselect2
	wire   [31:0] mm_interconnect_2_onchip_memory_s2_readdata;                                  // onchip_memory:readdata2 -> mm_interconnect_2:onchip_memory_s2_readdata
	wire   [15:0] mm_interconnect_2_onchip_memory_s2_address;                                   // mm_interconnect_2:onchip_memory_s2_address -> onchip_memory:address2
	wire    [3:0] mm_interconnect_2_onchip_memory_s2_byteenable;                                // mm_interconnect_2:onchip_memory_s2_byteenable -> onchip_memory:byteenable2
	wire          mm_interconnect_2_onchip_memory_s2_write;                                     // mm_interconnect_2:onchip_memory_s2_write -> onchip_memory:write2
	wire   [31:0] mm_interconnect_2_onchip_memory_s2_writedata;                                 // mm_interconnect_2:onchip_memory_s2_writedata -> onchip_memory:writedata2
	wire          mm_interconnect_2_onchip_memory_s2_clken;                                     // mm_interconnect_2:onchip_memory_s2_clken -> onchip_memory:clken2
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                              // hps_0:h2f_lw_AWBURST -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                                // hps_0:h2f_lw_ARLEN -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                                // hps_0:h2f_lw_WSTRB -> mm_interconnect_3:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                                               // mm_interconnect_3:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                                  // mm_interconnect_3:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                                               // hps_0:h2f_lw_RREADY -> mm_interconnect_3:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                                // hps_0:h2f_lw_AWLEN -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                                  // hps_0:h2f_lw_WID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                              // hps_0:h2f_lw_ARCACHE -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                                               // hps_0:h2f_lw_WVALID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                               // hps_0:h2f_lw_ARADDR -> mm_interconnect_3:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                               // hps_0:h2f_lw_ARPROT -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                               // hps_0:h2f_lw_AWPROT -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                                // hps_0:h2f_lw_WDATA -> mm_interconnect_3:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                                              // hps_0:h2f_lw_ARVALID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                              // hps_0:h2f_lw_AWCACHE -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                                 // hps_0:h2f_lw_ARID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                               // hps_0:h2f_lw_ARLOCK -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                               // hps_0:h2f_lw_AWLOCK -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                               // hps_0:h2f_lw_AWADDR -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                                // mm_interconnect_3:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                                              // mm_interconnect_3:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                                // mm_interconnect_3:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                                              // mm_interconnect_3:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                              // hps_0:h2f_lw_ARBURST -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                               // hps_0:h2f_lw_ARSIZE -> mm_interconnect_3:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                                               // hps_0:h2f_lw_BREADY -> mm_interconnect_3:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                                                // mm_interconnect_3:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                                                // hps_0:h2f_lw_WLAST -> mm_interconnect_3:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                                // mm_interconnect_3:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                                 // hps_0:h2f_lw_AWID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                                  // mm_interconnect_3:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                                               // mm_interconnect_3:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                               // hps_0:h2f_lw_AWSIZE -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                                              // hps_0:h2f_lw_AWVALID -> mm_interconnect_3:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                                               // mm_interconnect_3:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] master_non_sec_master_readdata;                                               // mm_interconnect_3:master_non_sec_master_readdata -> master_non_sec:master_readdata
	wire          master_non_sec_master_waitrequest;                                            // mm_interconnect_3:master_non_sec_master_waitrequest -> master_non_sec:master_waitrequest
	wire   [31:0] master_non_sec_master_address;                                                // master_non_sec:master_address -> mm_interconnect_3:master_non_sec_master_address
	wire          master_non_sec_master_read;                                                   // master_non_sec:master_read -> mm_interconnect_3:master_non_sec_master_read
	wire    [3:0] master_non_sec_master_byteenable;                                             // master_non_sec:master_byteenable -> mm_interconnect_3:master_non_sec_master_byteenable
	wire          master_non_sec_master_readdatavalid;                                          // mm_interconnect_3:master_non_sec_master_readdatavalid -> master_non_sec:master_readdatavalid
	wire          master_non_sec_master_write;                                                  // master_non_sec:master_write -> mm_interconnect_3:master_non_sec_master_write
	wire   [31:0] master_non_sec_master_writedata;                                              // master_non_sec:master_writedata -> mm_interconnect_3:master_non_sec_master_writedata
	wire   [31:0] mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_readdata;   // video_dma_controller_0:slave_readdata -> mm_interconnect_3:video_dma_controller_0_avalon_dma_control_slave_readdata
	wire    [1:0] mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_address;    // mm_interconnect_3:video_dma_controller_0_avalon_dma_control_slave_address -> video_dma_controller_0:slave_address
	wire          mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_read;       // mm_interconnect_3:video_dma_controller_0_avalon_dma_control_slave_read -> video_dma_controller_0:slave_read
	wire    [3:0] mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_byteenable; // mm_interconnect_3:video_dma_controller_0_avalon_dma_control_slave_byteenable -> video_dma_controller_0:slave_byteenable
	wire          mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_write;      // mm_interconnect_3:video_dma_controller_0_avalon_dma_control_slave_write -> video_dma_controller_0:slave_write
	wire   [31:0] mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_writedata;  // mm_interconnect_3:video_dma_controller_0_avalon_dma_control_slave_writedata -> video_dma_controller_0:slave_writedata
	wire          mm_interconnect_3_jtag_uart_avalon_jtag_slave_chipselect;                     // mm_interconnect_3:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_3_jtag_uart_avalon_jtag_slave_readdata;                       // jtag_uart:av_readdata -> mm_interconnect_3:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_3_jtag_uart_avalon_jtag_slave_waitrequest;                    // jtag_uart:av_waitrequest -> mm_interconnect_3:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_3_jtag_uart_avalon_jtag_slave_address;                        // mm_interconnect_3:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_3_jtag_uart_avalon_jtag_slave_read;                           // mm_interconnect_3:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_3_jtag_uart_avalon_jtag_slave_write;                          // mm_interconnect_3:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_3_jtag_uart_avalon_jtag_slave_writedata;                      // mm_interconnect_3:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [31:0] mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_readdata;                      // alt_vip_vfr_vga:slave_readdata -> mm_interconnect_3:alt_vip_vfr_vga_avalon_slave_readdata
	wire    [4:0] mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_address;                       // mm_interconnect_3:alt_vip_vfr_vga_avalon_slave_address -> alt_vip_vfr_vga:slave_address
	wire          mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_read;                          // mm_interconnect_3:alt_vip_vfr_vga_avalon_slave_read -> alt_vip_vfr_vga:slave_read
	wire          mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_write;                         // mm_interconnect_3:alt_vip_vfr_vga_avalon_slave_write -> alt_vip_vfr_vga:slave_write
	wire   [31:0] mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_writedata;                     // mm_interconnect_3:alt_vip_vfr_vga_avalon_slave_writedata -> alt_vip_vfr_vga:slave_writedata
	wire          mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_chipselect;               // mm_interconnect_3:i2c_opencores_mipi_avalon_slave_0_chipselect -> i2c_opencores_mipi:wb_stb_i
	wire    [7:0] mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_readdata;                 // i2c_opencores_mipi:wb_dat_o -> mm_interconnect_3:i2c_opencores_mipi_avalon_slave_0_readdata
	wire          mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_waitrequest;              // i2c_opencores_mipi:wb_ack_o -> mm_interconnect_3:i2c_opencores_mipi_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_address;                  // mm_interconnect_3:i2c_opencores_mipi_avalon_slave_0_address -> i2c_opencores_mipi:wb_adr_i
	wire          mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_write;                    // mm_interconnect_3:i2c_opencores_mipi_avalon_slave_0_write -> i2c_opencores_mipi:wb_we_i
	wire    [7:0] mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_writedata;                // mm_interconnect_3:i2c_opencores_mipi_avalon_slave_0_writedata -> i2c_opencores_mipi:wb_dat_i
	wire          mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_chipselect;             // mm_interconnect_3:i2c_opencores_camera_avalon_slave_0_chipselect -> i2c_opencores_camera:wb_stb_i
	wire    [7:0] mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_readdata;               // i2c_opencores_camera:wb_dat_o -> mm_interconnect_3:i2c_opencores_camera_avalon_slave_0_readdata
	wire          mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_waitrequest;            // i2c_opencores_camera:wb_ack_o -> mm_interconnect_3:i2c_opencores_camera_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_address;                // mm_interconnect_3:i2c_opencores_camera_avalon_slave_0_address -> i2c_opencores_camera:wb_adr_i
	wire          mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_write;                  // mm_interconnect_3:i2c_opencores_camera_avalon_slave_0_write -> i2c_opencores_camera:wb_we_i
	wire    [7:0] mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_writedata;              // mm_interconnect_3:i2c_opencores_camera_avalon_slave_0_writedata -> i2c_opencores_camera:wb_dat_i
	wire          mm_interconnect_3_alt_vip_mix_0_control_chipselect;                           // mm_interconnect_3:alt_vip_mix_0_control_chipselect -> alt_vip_mix_0:control_av_chipselect
	wire   [15:0] mm_interconnect_3_alt_vip_mix_0_control_readdata;                             // alt_vip_mix_0:control_av_readdata -> mm_interconnect_3:alt_vip_mix_0_control_readdata
	wire    [5:0] mm_interconnect_3_alt_vip_mix_0_control_address;                              // mm_interconnect_3:alt_vip_mix_0_control_address -> alt_vip_mix_0:control_av_address
	wire          mm_interconnect_3_alt_vip_mix_0_control_write;                                // mm_interconnect_3:alt_vip_mix_0_control_write -> alt_vip_mix_0:control_av_write
	wire   [15:0] mm_interconnect_3_alt_vip_mix_0_control_writedata;                            // mm_interconnect_3:alt_vip_mix_0_control_writedata -> alt_vip_mix_0:control_av_writedata
	wire   [31:0] mm_interconnect_3_alt_vip_cl_clp_1_control_readdata;                          // alt_vip_cl_clp_1:control_readdata -> mm_interconnect_3:alt_vip_cl_clp_1_control_readdata
	wire          mm_interconnect_3_alt_vip_cl_clp_1_control_waitrequest;                       // alt_vip_cl_clp_1:control_waitrequest -> mm_interconnect_3:alt_vip_cl_clp_1_control_waitrequest
	wire    [2:0] mm_interconnect_3_alt_vip_cl_clp_1_control_address;                           // mm_interconnect_3:alt_vip_cl_clp_1_control_address -> alt_vip_cl_clp_1:control_address
	wire          mm_interconnect_3_alt_vip_cl_clp_1_control_read;                              // mm_interconnect_3:alt_vip_cl_clp_1_control_read -> alt_vip_cl_clp_1:control_read
	wire    [3:0] mm_interconnect_3_alt_vip_cl_clp_1_control_byteenable;                        // mm_interconnect_3:alt_vip_cl_clp_1_control_byteenable -> alt_vip_cl_clp_1:control_byteenable
	wire          mm_interconnect_3_alt_vip_cl_clp_1_control_readdatavalid;                     // alt_vip_cl_clp_1:control_readdatavalid -> mm_interconnect_3:alt_vip_cl_clp_1_control_readdatavalid
	wire          mm_interconnect_3_alt_vip_cl_clp_1_control_write;                             // mm_interconnect_3:alt_vip_cl_clp_1_control_write -> alt_vip_cl_clp_1:control_write
	wire   [31:0] mm_interconnect_3_alt_vip_cl_clp_1_control_writedata;                         // mm_interconnect_3:alt_vip_cl_clp_1_control_writedata -> alt_vip_cl_clp_1:control_writedata
	wire   [31:0] mm_interconnect_3_sysid_qsys_control_slave_readdata;                          // sysid_qsys:readdata -> mm_interconnect_3:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_3_sysid_qsys_control_slave_address;                           // mm_interconnect_3:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire          mm_interconnect_3_led_s1_chipselect;                                          // mm_interconnect_3:led_s1_chipselect -> led:chipselect
	wire   [31:0] mm_interconnect_3_led_s1_readdata;                                            // led:readdata -> mm_interconnect_3:led_s1_readdata
	wire    [1:0] mm_interconnect_3_led_s1_address;                                             // mm_interconnect_3:led_s1_address -> led:address
	wire          mm_interconnect_3_led_s1_write;                                               // mm_interconnect_3:led_s1_write -> led:write_n
	wire   [31:0] mm_interconnect_3_led_s1_writedata;                                           // mm_interconnect_3:led_s1_writedata -> led:writedata
	wire          mm_interconnect_3_sw_s1_chipselect;                                           // mm_interconnect_3:sw_s1_chipselect -> sw:chipselect
	wire   [31:0] mm_interconnect_3_sw_s1_readdata;                                             // sw:readdata -> mm_interconnect_3:sw_s1_readdata
	wire    [1:0] mm_interconnect_3_sw_s1_address;                                              // mm_interconnect_3:sw_s1_address -> sw:address
	wire          mm_interconnect_3_sw_s1_write;                                                // mm_interconnect_3:sw_s1_write -> sw:write_n
	wire   [31:0] mm_interconnect_3_sw_s1_writedata;                                            // mm_interconnect_3:sw_s1_writedata -> sw:writedata
	wire          mm_interconnect_3_key_s1_chipselect;                                          // mm_interconnect_3:key_s1_chipselect -> key:chipselect
	wire   [31:0] mm_interconnect_3_key_s1_readdata;                                            // key:readdata -> mm_interconnect_3:key_s1_readdata
	wire    [1:0] mm_interconnect_3_key_s1_address;                                             // mm_interconnect_3:key_s1_address -> key:address
	wire          mm_interconnect_3_key_s1_write;                                               // mm_interconnect_3:key_s1_write -> key:write_n
	wire   [31:0] mm_interconnect_3_key_s1_writedata;                                           // mm_interconnect_3:key_s1_writedata -> key:writedata
	wire          mm_interconnect_3_mipi_reset_n_s1_chipselect;                                 // mm_interconnect_3:mipi_reset_n_s1_chipselect -> mipi_reset_n:chipselect
	wire   [31:0] mm_interconnect_3_mipi_reset_n_s1_readdata;                                   // mipi_reset_n:readdata -> mm_interconnect_3:mipi_reset_n_s1_readdata
	wire    [1:0] mm_interconnect_3_mipi_reset_n_s1_address;                                    // mm_interconnect_3:mipi_reset_n_s1_address -> mipi_reset_n:address
	wire          mm_interconnect_3_mipi_reset_n_s1_write;                                      // mm_interconnect_3:mipi_reset_n_s1_write -> mipi_reset_n:write_n
	wire   [31:0] mm_interconnect_3_mipi_reset_n_s1_writedata;                                  // mm_interconnect_3:mipi_reset_n_s1_writedata -> mipi_reset_n:writedata
	wire          mm_interconnect_3_mipi_pwdn_n_s1_chipselect;                                  // mm_interconnect_3:mipi_pwdn_n_s1_chipselect -> mipi_pwdn_n:chipselect
	wire   [31:0] mm_interconnect_3_mipi_pwdn_n_s1_readdata;                                    // mipi_pwdn_n:readdata -> mm_interconnect_3:mipi_pwdn_n_s1_readdata
	wire    [1:0] mm_interconnect_3_mipi_pwdn_n_s1_address;                                     // mm_interconnect_3:mipi_pwdn_n_s1_address -> mipi_pwdn_n:address
	wire          mm_interconnect_3_mipi_pwdn_n_s1_write;                                       // mm_interconnect_3:mipi_pwdn_n_s1_write -> mipi_pwdn_n:write_n
	wire   [31:0] mm_interconnect_3_mipi_pwdn_n_s1_writedata;                                   // mm_interconnect_3:mipi_pwdn_n_s1_writedata -> mipi_pwdn_n:writedata
	wire   [31:0] mm_interconnect_3_intr_capturer_0_avalon_slave_0_readdata;                    // intr_capturer_0:rddata -> mm_interconnect_3:intr_capturer_0_avalon_slave_0_readdata
	wire    [0:0] mm_interconnect_3_intr_capturer_0_avalon_slave_0_address;                     // mm_interconnect_3:intr_capturer_0_avalon_slave_0_address -> intr_capturer_0:addr
	wire          mm_interconnect_3_intr_capturer_0_avalon_slave_0_read;                        // mm_interconnect_3:intr_capturer_0_avalon_slave_0_read -> intr_capturer_0:read
	wire   [31:0] hps_0_f2h_irq0_irq;                                                           // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                                           // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire   [31:0] intr_capturer_0_interrupt_receiver_irq;                                       // irq_mapper_002:sender_irq -> intr_capturer_0:interrupt_in
	wire          irq_mapper_receiver0_irq;                                                     // jtag_uart:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_002:receiver0_irq]
	wire          irq_mapper_receiver1_irq;                                                     // key:irq -> [irq_mapper:receiver1_irq, irq_mapper_002:receiver1_irq]
	wire          irq_mapper_receiver2_irq;                                                     // sw:irq -> [irq_mapper:receiver2_irq, irq_mapper_002:receiver2_irq]
	wire          rst_controller_reset_out_reset;                                               // rst_controller:reset_out -> [TERASIC_CAMERA_0:reset_n, alt_vip_cl_clp_1:main_reset, alt_vip_cl_scl_0:main_reset, alt_vip_cl_tpg_0:main_reset, alt_vip_cpr_0:reset, alt_vip_cpr_1:reset, alt_vip_cpr_2:reset, alt_vip_itc_0:rst, alt_vip_mix_0:reset, alt_vip_vfb_0:reset, alt_vip_vfr_vga:master_reset, alt_vip_vfr_vga:reset, mm_interconnect_0:video_dma_controller_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset_reset, mm_interconnect_2:alt_vip_vfb_0_reset_reset_bridge_in_reset_reset, mm_interconnect_3:video_dma_controller_0_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_translator:in_reset, sdram:reset_n, st_adapter_0:in_rst_0_reset, video_csc_0:reset, video_dma_controller_0:reset]
	wire          rst_controller_reset_out_reset_req;                                           // rst_controller:reset_req -> [onchip_memory:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                                           // rst_controller_001:reset_out -> [i2c_opencores_camera:wb_rst_i, i2c_opencores_mipi:wb_rst_i, intr_capturer_0:rst_n, irq_mapper_002:reset, jtag_uart:rst_n, key:reset_n, led:reset_n, mipi_pwdn_n:reset_n, mipi_reset_n:reset_n, mm_interconnect_1:master_secure_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:master_secure_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_3:jtag_uart_reset_reset_bridge_in_reset_reset, mm_interconnect_3:master_non_sec_clk_reset_reset_bridge_in_reset_reset, sw:reset_n, sysid_qsys:reset_n]
	wire          rst_controller_002_reset_out_reset;                                           // rst_controller_002:reset_out -> [mm_interconnect_1:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_3:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	TERASIC_CAMERA #(
		.VIDEO_W (640),
		.VIDEO_H (480)
	) terasic_camera_0 (
		.clk           (pll_0_outclk0_clk),                                      //             clock_reset.clk
		.reset_n       (~rst_controller_reset_out_reset),                        //       clock_reset_reset.reset_n
		.CAMERA_D      (terasic_camera_0_conduit_end_D),                         //             conduit_end.export
		.CAMERA_FVAL   (terasic_camera_0_conduit_end_FVAL),                      //                        .export
		.CAMERA_LVAL   (terasic_camera_0_conduit_end_LVAL),                      //                        .export
		.CAMERA_PIXCLK (terasic_camera_0_conduit_end_PIXCLK),                    //                        .export
		.st_data       (terasic_camera_0_avalon_streaming_source_data),          // avalon_streaming_source.data
		.st_sop        (terasic_camera_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.st_eop        (terasic_camera_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.st_ready      (terasic_camera_0_avalon_streaming_source_ready),         //                        .ready
		.st_valid      (terasic_camera_0_avalon_streaming_source_valid)          //                        .valid
	);

	soc_system_alt_vip_cl_clp_1 #(
		.MAX_IN_WIDTH                 (640),
		.MAX_IN_HEIGHT                (480),
		.BITS_PER_SYMBOL              (8),
		.PIXELS_IN_PARALLEL           (1),
		.NUMBER_OF_COLOR_PLANES       (3),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.CLIPPING_METHOD              ("RECTANGLE"),
		.LEFT_OFFSET                  (0),
		.RIGHT_OFFSET                 (10),
		.TOP_OFFSET                   (0),
		.BOTTOM_OFFSET                (10),
		.RECTANGLE_WIDTH              (640),
		.RECTANGLE_HEIGHT             (480),
		.RUNTIME_CONTROL              (1)
	) alt_vip_cl_clp_1 (
		.main_clock            (pll_0_outclk0_clk),                                        // main_clock.clk
		.main_reset            (rst_controller_reset_out_reset),                           // main_reset.reset
		.din_data              (terasic_camera_0_avalon_streaming_source_data),            //        din.data
		.din_valid             (terasic_camera_0_avalon_streaming_source_valid),           //           .valid
		.din_startofpacket     (terasic_camera_0_avalon_streaming_source_startofpacket),   //           .startofpacket
		.din_endofpacket       (terasic_camera_0_avalon_streaming_source_endofpacket),     //           .endofpacket
		.din_ready             (terasic_camera_0_avalon_streaming_source_ready),           //           .ready
		.dout_data             (alt_vip_cl_clp_1_dout_data),                               //       dout.data
		.dout_valid            (alt_vip_cl_clp_1_dout_valid),                              //           .valid
		.dout_startofpacket    (alt_vip_cl_clp_1_dout_startofpacket),                      //           .startofpacket
		.dout_endofpacket      (alt_vip_cl_clp_1_dout_endofpacket),                        //           .endofpacket
		.dout_ready            (alt_vip_cl_clp_1_dout_ready),                              //           .ready
		.control_address       (mm_interconnect_3_alt_vip_cl_clp_1_control_address),       //    control.address
		.control_byteenable    (mm_interconnect_3_alt_vip_cl_clp_1_control_byteenable),    //           .byteenable
		.control_write         (mm_interconnect_3_alt_vip_cl_clp_1_control_write),         //           .write
		.control_writedata     (mm_interconnect_3_alt_vip_cl_clp_1_control_writedata),     //           .writedata
		.control_read          (mm_interconnect_3_alt_vip_cl_clp_1_control_read),          //           .read
		.control_readdata      (mm_interconnect_3_alt_vip_cl_clp_1_control_readdata),      //           .readdata
		.control_readdatavalid (mm_interconnect_3_alt_vip_cl_clp_1_control_readdatavalid), //           .readdatavalid
		.control_waitrequest   (mm_interconnect_3_alt_vip_cl_clp_1_control_waitrequest)    //           .waitrequest
	);

	soc_system_alt_vip_cl_scl_0 #(
		.SYMBOLS_IN_SEQ      (1),
		.SYMBOLS_IN_PAR      (3),
		.BITS_PER_SYMBOL     (8),
		.EXTRA_PIPELINING    (0),
		.IS_422              (1),
		.NO_BLANKING         (0),
		.MAX_IN_WIDTH        (640),
		.MAX_IN_HEIGHT       (480),
		.MAX_OUT_WIDTH       (320),
		.MAX_OUT_HEIGHT      (240),
		.RUNTIME_CONTROL     (0),
		.ALWAYS_DOWNSCALE    (0),
		.ALGORITHM_NAME      ("POLYPHASE"),
		.DEFAULT_EDGE_THRESH (7),
		.DEFAULT_UPPER_BLUR  (15),
		.DEFAULT_LOWER_BLUR  (0),
		.ENABLE_FIR          (0),
		.ARE_IDENTICAL       (0),
		.V_TAPS              (8),
		.V_PHASES            (16),
		.H_TAPS              (8),
		.H_PHASES            (16),
		.V_SIGNED            (1),
		.V_INTEGER_BITS      (1),
		.V_FRACTION_BITS     (7),
		.H_SIGNED            (1),
		.H_INTEGER_BITS      (1),
		.H_FRACTION_BITS     (7),
		.PRESERVE_BITS       (0),
		.LOAD_AT_RUNTIME     (0),
		.V_BANKS             (1),
		.V_SYMMETRIC         (0),
		.V_FUNCTION          ("LANCZOS_2"),
		.V_COEFF_FILE        ("<enter file name (including full path)>"),
		.H_BANKS             (1),
		.H_SYMMETRIC         (0),
		.H_FUNCTION          ("LANCZOS_2"),
		.H_COEFF_FILE        ("<enter file name (including full path)>"),
		.IS_420              (0)
	) alt_vip_cl_scl_0 (
		.main_clock         (pll_0_outclk0_clk),                   // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.din_data           (alt_vip_cl_clp_1_dout_data),          //        din.data
		.din_valid          (alt_vip_cl_clp_1_dout_valid),         //           .valid
		.din_startofpacket  (alt_vip_cl_clp_1_dout_startofpacket), //           .startofpacket
		.din_endofpacket    (alt_vip_cl_clp_1_dout_endofpacket),   //           .endofpacket
		.din_ready          (alt_vip_cl_clp_1_dout_ready),         //           .ready
		.dout_data          (alt_vip_cl_scl_0_dout_data),          //       dout.data
		.dout_valid         (alt_vip_cl_scl_0_dout_valid),         //           .valid
		.dout_startofpacket (alt_vip_cl_scl_0_dout_startofpacket), //           .startofpacket
		.dout_endofpacket   (alt_vip_cl_scl_0_dout_endofpacket),   //           .endofpacket
		.dout_ready         (alt_vip_cl_scl_0_dout_ready)          //           .ready
	);

	soc_system_alt_vip_cl_tpg_0 #(
		.BPS                          (8),
		.PIXELS_IN_PARALLEL           (1),
		.MAX_WIDTH                    (640),
		.MAX_HEIGHT                   (480),
		.OUTPUT_FORMAT                ("4.4.4"),
		.COLOR_SPACE                  ("RGB"),
		.INTERLACING                  ("prog"),
		.PATTERN                      ("colorbars"),
		.UNIFORM_VALUE_RY             (16),
		.UNIFORM_VALUE_GCB            (16),
		.UNIFORM_VALUE_BCR            (16),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.RUNTIME_CONTROL              (0)
	) alt_vip_cl_tpg_0 (
		.main_clock         (pll_0_outclk0_clk),                   // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.dout_data          (alt_vip_cl_tpg_0_dout_data),          //       dout.data
		.dout_valid         (alt_vip_cl_tpg_0_dout_valid),         //           .valid
		.dout_startofpacket (alt_vip_cl_tpg_0_dout_startofpacket), //           .startofpacket
		.dout_endofpacket   (alt_vip_cl_tpg_0_dout_endofpacket),   //           .endofpacket
		.dout_ready         (alt_vip_cl_tpg_0_dout_ready)          //           .ready
	);

	soc_system_alt_vip_cpr_0 alt_vip_cpr_0 (
		.clock               (pll_0_outclk0_clk),                                     // clock.clk
		.reset               (rst_controller_reset_out_reset),                        // reset.reset
		.din0_ready          (alt_vip_vfr_vga_avalon_streaming_source_ready),         //  din0.ready
		.din0_valid          (alt_vip_vfr_vga_avalon_streaming_source_valid),         //      .valid
		.din0_data           (alt_vip_vfr_vga_avalon_streaming_source_data),          //      .data
		.din0_startofpacket  (alt_vip_vfr_vga_avalon_streaming_source_startofpacket), //      .startofpacket
		.din0_endofpacket    (alt_vip_vfr_vga_avalon_streaming_source_endofpacket),   //      .endofpacket
		.dout0_ready         (alt_vip_cpr_0_dout0_ready),                             // dout0.ready
		.dout0_valid         (alt_vip_cpr_0_dout0_valid),                             //      .valid
		.dout0_data          (alt_vip_cpr_0_dout0_data),                              //      .data
		.dout0_startofpacket (alt_vip_cpr_0_dout0_startofpacket),                     //      .startofpacket
		.dout0_endofpacket   (alt_vip_cpr_0_dout0_endofpacket)                        //      .endofpacket
	);

	soc_system_alt_vip_cpr_1 alt_vip_cpr_1 (
		.clock               (pll_0_outclk0_clk),                 // clock.clk
		.reset               (rst_controller_reset_out_reset),    // reset.reset
		.din0_ready          (alt_vip_cpr_2_dout0_ready),         //  din0.ready
		.din0_valid          (alt_vip_cpr_2_dout0_valid),         //      .valid
		.din0_data           (alt_vip_cpr_2_dout0_data),          //      .data
		.din0_startofpacket  (alt_vip_cpr_2_dout0_startofpacket), //      .startofpacket
		.din0_endofpacket    (alt_vip_cpr_2_dout0_endofpacket),   //      .endofpacket
		.dout0_ready         (alt_vip_cpr_1_dout0_ready),         // dout0.ready
		.dout0_valid         (alt_vip_cpr_1_dout0_valid),         //      .valid
		.dout0_data          (alt_vip_cpr_1_dout0_data),          //      .data
		.dout0_startofpacket (alt_vip_cpr_1_dout0_startofpacket), //      .startofpacket
		.dout0_endofpacket   (alt_vip_cpr_1_dout0_endofpacket)    //      .endofpacket
	);

	soc_system_alt_vip_cpr_2 alt_vip_cpr_2 (
		.clock               (pll_0_outclk0_clk),                 // clock.clk
		.reset               (rst_controller_reset_out_reset),    // reset.reset
		.din0_ready          (alt_vip_vfb_0_dout_ready),          //  din0.ready
		.din0_valid          (alt_vip_vfb_0_dout_valid),          //      .valid
		.din0_data           (alt_vip_vfb_0_dout_data),           //      .data
		.din0_startofpacket  (alt_vip_vfb_0_dout_startofpacket),  //      .startofpacket
		.din0_endofpacket    (alt_vip_vfb_0_dout_endofpacket),    //      .endofpacket
		.dout0_ready         (alt_vip_cpr_2_dout0_ready),         // dout0.ready
		.dout0_valid         (alt_vip_cpr_2_dout0_valid),         //      .valid
		.dout0_data          (alt_vip_cpr_2_dout0_data),          //      .data
		.dout0_startofpacket (alt_vip_cpr_2_dout0_startofpacket), //      .startofpacket
		.dout0_endofpacket   (alt_vip_cpr_2_dout0_endofpacket),   //      .endofpacket
		.dout1_ready         (alt_vip_cpr_2_dout1_ready),         // dout1.ready
		.dout1_valid         (alt_vip_cpr_2_dout1_valid),         //      .valid
		.dout1_data          (alt_vip_cpr_2_dout1_data),          //      .data
		.dout1_startofpacket (alt_vip_cpr_2_dout1_startofpacket), //      .startofpacket
		.dout1_endofpacket   (alt_vip_cpr_2_dout1_endofpacket)    //      .endofpacket
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (1024),
		.V_ACTIVE_LINES                (768),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (10240),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (10239),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (136),
		.H_FRONT_PORCH                 (24),
		.H_BACK_PORCH                  (160),
		.V_SYNC_LENGTH                 (6),
		.V_FRONT_PORCH                 (3),
		.V_BACK_PORCH                  (29),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (pll_0_outclk0_clk),                         //       is_clk_rst.clk
		.rst           (rst_controller_reset_out_reset),            // is_clk_rst_reset.reset
		.is_data       (alt_vip_mix_0_dout_data),                   //              din.data
		.is_valid      (alt_vip_mix_0_dout_valid),                  //                 .valid
		.is_ready      (alt_vip_mix_0_dout_ready),                  //                 .ready
		.is_sop        (alt_vip_mix_0_dout_startofpacket),          //                 .startofpacket
		.is_eop        (alt_vip_mix_0_dout_endofpacket),            //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),       //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),      //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),     //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid), //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),    //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),    //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),         //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),         //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)          //                 .export
	);

	soc_system_alt_vip_mix_0 alt_vip_mix_0 (
		.clock                 (pll_0_outclk0_clk),                                  //   clock.clk
		.reset                 (rst_controller_reset_out_reset),                     //   reset.reset
		.din_0_ready           (alt_vip_cpr_0_dout0_ready),                          //   din_0.ready
		.din_0_valid           (alt_vip_cpr_0_dout0_valid),                          //        .valid
		.din_0_data            (alt_vip_cpr_0_dout0_data),                           //        .data
		.din_0_startofpacket   (alt_vip_cpr_0_dout0_startofpacket),                  //        .startofpacket
		.din_0_endofpacket     (alt_vip_cpr_0_dout0_endofpacket),                    //        .endofpacket
		.din_1_ready           (alt_vip_cpr_1_dout0_ready),                          //   din_1.ready
		.din_1_valid           (alt_vip_cpr_1_dout0_valid),                          //        .valid
		.din_1_data            (alt_vip_cpr_1_dout0_data),                           //        .data
		.din_1_startofpacket   (alt_vip_cpr_1_dout0_startofpacket),                  //        .startofpacket
		.din_1_endofpacket     (alt_vip_cpr_1_dout0_endofpacket),                    //        .endofpacket
		.din_2_ready           (alt_vip_cl_tpg_0_dout_ready),                        //   din_2.ready
		.din_2_valid           (alt_vip_cl_tpg_0_dout_valid),                        //        .valid
		.din_2_data            (alt_vip_cl_tpg_0_dout_data),                         //        .data
		.din_2_startofpacket   (alt_vip_cl_tpg_0_dout_startofpacket),                //        .startofpacket
		.din_2_endofpacket     (alt_vip_cl_tpg_0_dout_endofpacket),                  //        .endofpacket
		.dout_ready            (alt_vip_mix_0_dout_ready),                           //    dout.ready
		.dout_valid            (alt_vip_mix_0_dout_valid),                           //        .valid
		.dout_data             (alt_vip_mix_0_dout_data),                            //        .data
		.dout_startofpacket    (alt_vip_mix_0_dout_startofpacket),                   //        .startofpacket
		.dout_endofpacket      (alt_vip_mix_0_dout_endofpacket),                     //        .endofpacket
		.control_av_chipselect (mm_interconnect_3_alt_vip_mix_0_control_chipselect), // control.chipselect
		.control_av_write      (mm_interconnect_3_alt_vip_mix_0_control_write),      //        .write
		.control_av_address    (mm_interconnect_3_alt_vip_mix_0_control_address),    //        .address
		.control_av_writedata  (mm_interconnect_3_alt_vip_mix_0_control_writedata),  //        .writedata
		.control_av_readdata   (mm_interconnect_3_alt_vip_mix_0_control_readdata)    //        .readdata
	);

	soc_system_alt_vip_vfb_0 alt_vip_vfb_0 (
		.clock                        (pll_0_outclk0_clk),                       //        clock.clk
		.reset                        (rst_controller_reset_out_reset),          //        reset.reset
		.din_ready                    (alt_vip_cl_scl_0_dout_ready),             //          din.ready
		.din_valid                    (alt_vip_cl_scl_0_dout_valid),             //             .valid
		.din_data                     (alt_vip_cl_scl_0_dout_data),              //             .data
		.din_startofpacket            (alt_vip_cl_scl_0_dout_startofpacket),     //             .startofpacket
		.din_endofpacket              (alt_vip_cl_scl_0_dout_endofpacket),       //             .endofpacket
		.dout_ready                   (alt_vip_vfb_0_dout_ready),                //         dout.ready
		.dout_valid                   (alt_vip_vfb_0_dout_valid),                //             .valid
		.dout_data                    (alt_vip_vfb_0_dout_data),                 //             .data
		.dout_startofpacket           (alt_vip_vfb_0_dout_startofpacket),        //             .startofpacket
		.dout_endofpacket             (alt_vip_vfb_0_dout_endofpacket),          //             .endofpacket
		.read_master_av_address       (alt_vip_vfb_0_read_master_address),       //  read_master.address
		.read_master_av_read          (alt_vip_vfb_0_read_master_read),          //             .read
		.read_master_av_waitrequest   (alt_vip_vfb_0_read_master_waitrequest),   //             .waitrequest
		.read_master_av_readdatavalid (alt_vip_vfb_0_read_master_readdatavalid), //             .readdatavalid
		.read_master_av_readdata      (alt_vip_vfb_0_read_master_readdata),      //             .readdata
		.read_master_av_burstcount    (alt_vip_vfb_0_read_master_burstcount),    //             .burstcount
		.write_master_av_address      (alt_vip_vfb_0_write_master_address),      // write_master.address
		.write_master_av_write        (alt_vip_vfb_0_write_master_write),        //             .write
		.write_master_av_writedata    (alt_vip_vfb_0_write_master_writedata),    //             .writedata
		.write_master_av_waitrequest  (alt_vip_vfb_0_write_master_waitrequest),  //             .waitrequest
		.write_master_av_burstcount   (alt_vip_vfb_0_write_master_burstcount)    //             .burstcount
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (4),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (1024),
		.MAX_IMAGE_HEIGHT               (768),
		.MEM_PORT_WIDTH                 (128),
		.RMASTER_FIFO_DEPTH             (64),
		.RMASTER_BURST_TARGET           (32),
		.CLOCKS_ARE_SEPARATE            (1)
	) alt_vip_vfr_vga (
		.clock                (pll_0_outclk0_clk),                                        //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                           //       clock_reset_reset.reset
		.master_clock         (pll_0_outclk0_clk),                                        //            clock_master.clk
		.master_reset         (rst_controller_reset_out_reset),                           //      clock_master_reset.reset
		.slave_address        (mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (),                                                         //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_vga_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_vga_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_vga_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_vga_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_vga_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_vga_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_vga_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_vga_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_vga_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_vga_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_vga_avalon_master_waitrequest)                 //                        .waitrequest
	);

	soc_system_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (2)
	) hps_0 (
		.f2h_boot_from_fpga_ready      (),                                              // f2h_boot_from_fpga.boot_from_fpga_ready
		.f2h_boot_from_fpga_on_failure (),                                              //                   .boot_from_fpga_on_failure
		.mem_a                         (memory_mem_a),                                  //             memory.mem_a
		.mem_ba                        (memory_mem_ba),                                 //                   .mem_ba
		.mem_ck                        (memory_mem_ck),                                 //                   .mem_ck
		.mem_ck_n                      (memory_mem_ck_n),                               //                   .mem_ck_n
		.mem_cke                       (memory_mem_cke),                                //                   .mem_cke
		.mem_cs_n                      (memory_mem_cs_n),                               //                   .mem_cs_n
		.mem_ras_n                     (memory_mem_ras_n),                              //                   .mem_ras_n
		.mem_cas_n                     (memory_mem_cas_n),                              //                   .mem_cas_n
		.mem_we_n                      (memory_mem_we_n),                               //                   .mem_we_n
		.mem_reset_n                   (memory_mem_reset_n),                            //                   .mem_reset_n
		.mem_dq                        (memory_mem_dq),                                 //                   .mem_dq
		.mem_dqs                       (memory_mem_dqs),                                //                   .mem_dqs
		.mem_dqs_n                     (memory_mem_dqs_n),                              //                   .mem_dqs_n
		.mem_odt                       (memory_mem_odt),                                //                   .mem_odt
		.mem_dm                        (memory_mem_dm),                                 //                   .mem_dm
		.oct_rzqin                     (memory_oct_rzqin),                              //                   .oct_rzqin
		.hps_io_emac1_inst_TX_CLK      (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),         //             hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0        (hps_0_hps_io_hps_io_emac1_inst_TXD0),           //                   .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1        (hps_0_hps_io_hps_io_emac1_inst_TXD1),           //                   .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2        (hps_0_hps_io_hps_io_emac1_inst_TXD2),           //                   .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3        (hps_0_hps_io_hps_io_emac1_inst_TXD3),           //                   .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0        (hps_0_hps_io_hps_io_emac1_inst_RXD0),           //                   .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO        (hps_0_hps_io_hps_io_emac1_inst_MDIO),           //                   .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC         (hps_0_hps_io_hps_io_emac1_inst_MDC),            //                   .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL      (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),         //                   .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL      (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),         //                   .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK      (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),         //                   .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1        (hps_0_hps_io_hps_io_emac1_inst_RXD1),           //                   .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2        (hps_0_hps_io_hps_io_emac1_inst_RXD2),           //                   .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3        (hps_0_hps_io_hps_io_emac1_inst_RXD3),           //                   .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0          (hps_0_hps_io_hps_io_qspi_inst_IO0),             //                   .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1          (hps_0_hps_io_hps_io_qspi_inst_IO1),             //                   .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2          (hps_0_hps_io_hps_io_qspi_inst_IO2),             //                   .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3          (hps_0_hps_io_hps_io_qspi_inst_IO3),             //                   .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0          (hps_0_hps_io_hps_io_qspi_inst_SS0),             //                   .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK          (hps_0_hps_io_hps_io_qspi_inst_CLK),             //                   .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD          (hps_0_hps_io_hps_io_sdio_inst_CMD),             //                   .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0           (hps_0_hps_io_hps_io_sdio_inst_D0),              //                   .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1           (hps_0_hps_io_hps_io_sdio_inst_D1),              //                   .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK          (hps_0_hps_io_hps_io_sdio_inst_CLK),             //                   .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2           (hps_0_hps_io_hps_io_sdio_inst_D2),              //                   .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3           (hps_0_hps_io_hps_io_sdio_inst_D3),              //                   .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0           (hps_0_hps_io_hps_io_usb1_inst_D0),              //                   .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1           (hps_0_hps_io_hps_io_usb1_inst_D1),              //                   .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2           (hps_0_hps_io_hps_io_usb1_inst_D2),              //                   .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3           (hps_0_hps_io_hps_io_usb1_inst_D3),              //                   .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4           (hps_0_hps_io_hps_io_usb1_inst_D4),              //                   .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5           (hps_0_hps_io_hps_io_usb1_inst_D5),              //                   .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6           (hps_0_hps_io_hps_io_usb1_inst_D6),              //                   .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7           (hps_0_hps_io_hps_io_usb1_inst_D7),              //                   .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK          (hps_0_hps_io_hps_io_usb1_inst_CLK),             //                   .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP          (hps_0_hps_io_hps_io_usb1_inst_STP),             //                   .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR          (hps_0_hps_io_hps_io_usb1_inst_DIR),             //                   .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT          (hps_0_hps_io_hps_io_usb1_inst_NXT),             //                   .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK         (hps_0_hps_io_hps_io_spim1_inst_CLK),            //                   .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI        (hps_0_hps_io_hps_io_spim1_inst_MOSI),           //                   .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO        (hps_0_hps_io_hps_io_spim1_inst_MISO),           //                   .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0         (hps_0_hps_io_hps_io_spim1_inst_SS0),            //                   .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX          (hps_0_hps_io_hps_io_uart0_inst_RX),             //                   .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX          (hps_0_hps_io_hps_io_uart0_inst_TX),             //                   .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA          (hps_0_hps_io_hps_io_i2c0_inst_SDA),             //                   .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL          (hps_0_hps_io_hps_io_i2c0_inst_SCL),             //                   .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA          (hps_0_hps_io_hps_io_i2c1_inst_SDA),             //                   .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL          (hps_0_hps_io_hps_io_i2c1_inst_SCL),             //                   .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09       (hps_0_hps_io_hps_io_gpio_inst_GPIO09),          //                   .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35       (hps_0_hps_io_hps_io_gpio_inst_GPIO35),          //                   .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40       (hps_0_hps_io_hps_io_gpio_inst_GPIO40),          //                   .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48       (hps_0_hps_io_hps_io_gpio_inst_GPIO48),          //                   .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53       (hps_0_hps_io_hps_io_gpio_inst_GPIO53),          //                   .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54       (hps_0_hps_io_hps_io_gpio_inst_GPIO54),          //                   .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61       (hps_0_hps_io_hps_io_gpio_inst_GPIO61),          //                   .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                     (hps_0_h2f_reset_reset_n),                       //          h2f_reset.reset_n
		.h2f_axi_clk                   (clk_clk),                                       //      h2f_axi_clock.clk
		.h2f_AWID                      (hps_0_h2f_axi_master_awid),                     //     h2f_axi_master.awid
		.h2f_AWADDR                    (hps_0_h2f_axi_master_awaddr),                   //                   .awaddr
		.h2f_AWLEN                     (hps_0_h2f_axi_master_awlen),                    //                   .awlen
		.h2f_AWSIZE                    (hps_0_h2f_axi_master_awsize),                   //                   .awsize
		.h2f_AWBURST                   (hps_0_h2f_axi_master_awburst),                  //                   .awburst
		.h2f_AWLOCK                    (hps_0_h2f_axi_master_awlock),                   //                   .awlock
		.h2f_AWCACHE                   (hps_0_h2f_axi_master_awcache),                  //                   .awcache
		.h2f_AWPROT                    (hps_0_h2f_axi_master_awprot),                   //                   .awprot
		.h2f_AWVALID                   (hps_0_h2f_axi_master_awvalid),                  //                   .awvalid
		.h2f_AWREADY                   (hps_0_h2f_axi_master_awready),                  //                   .awready
		.h2f_WID                       (hps_0_h2f_axi_master_wid),                      //                   .wid
		.h2f_WDATA                     (hps_0_h2f_axi_master_wdata),                    //                   .wdata
		.h2f_WSTRB                     (hps_0_h2f_axi_master_wstrb),                    //                   .wstrb
		.h2f_WLAST                     (hps_0_h2f_axi_master_wlast),                    //                   .wlast
		.h2f_WVALID                    (hps_0_h2f_axi_master_wvalid),                   //                   .wvalid
		.h2f_WREADY                    (hps_0_h2f_axi_master_wready),                   //                   .wready
		.h2f_BID                       (hps_0_h2f_axi_master_bid),                      //                   .bid
		.h2f_BRESP                     (hps_0_h2f_axi_master_bresp),                    //                   .bresp
		.h2f_BVALID                    (hps_0_h2f_axi_master_bvalid),                   //                   .bvalid
		.h2f_BREADY                    (hps_0_h2f_axi_master_bready),                   //                   .bready
		.h2f_ARID                      (hps_0_h2f_axi_master_arid),                     //                   .arid
		.h2f_ARADDR                    (hps_0_h2f_axi_master_araddr),                   //                   .araddr
		.h2f_ARLEN                     (hps_0_h2f_axi_master_arlen),                    //                   .arlen
		.h2f_ARSIZE                    (hps_0_h2f_axi_master_arsize),                   //                   .arsize
		.h2f_ARBURST                   (hps_0_h2f_axi_master_arburst),                  //                   .arburst
		.h2f_ARLOCK                    (hps_0_h2f_axi_master_arlock),                   //                   .arlock
		.h2f_ARCACHE                   (hps_0_h2f_axi_master_arcache),                  //                   .arcache
		.h2f_ARPROT                    (hps_0_h2f_axi_master_arprot),                   //                   .arprot
		.h2f_ARVALID                   (hps_0_h2f_axi_master_arvalid),                  //                   .arvalid
		.h2f_ARREADY                   (hps_0_h2f_axi_master_arready),                  //                   .arready
		.h2f_RID                       (hps_0_h2f_axi_master_rid),                      //                   .rid
		.h2f_RDATA                     (hps_0_h2f_axi_master_rdata),                    //                   .rdata
		.h2f_RRESP                     (hps_0_h2f_axi_master_rresp),                    //                   .rresp
		.h2f_RLAST                     (hps_0_h2f_axi_master_rlast),                    //                   .rlast
		.h2f_RVALID                    (hps_0_h2f_axi_master_rvalid),                   //                   .rvalid
		.h2f_RREADY                    (hps_0_h2f_axi_master_rready),                   //                   .rready
		.f2h_axi_clk                   (clk_clk),                                       //      f2h_axi_clock.clk
		.f2h_AWID                      (mm_interconnect_1_hps_0_f2h_axi_slave_awid),    //      f2h_axi_slave.awid
		.f2h_AWADDR                    (mm_interconnect_1_hps_0_f2h_axi_slave_awaddr),  //                   .awaddr
		.f2h_AWLEN                     (mm_interconnect_1_hps_0_f2h_axi_slave_awlen),   //                   .awlen
		.f2h_AWSIZE                    (mm_interconnect_1_hps_0_f2h_axi_slave_awsize),  //                   .awsize
		.f2h_AWBURST                   (mm_interconnect_1_hps_0_f2h_axi_slave_awburst), //                   .awburst
		.f2h_AWLOCK                    (mm_interconnect_1_hps_0_f2h_axi_slave_awlock),  //                   .awlock
		.f2h_AWCACHE                   (mm_interconnect_1_hps_0_f2h_axi_slave_awcache), //                   .awcache
		.f2h_AWPROT                    (mm_interconnect_1_hps_0_f2h_axi_slave_awprot),  //                   .awprot
		.f2h_AWVALID                   (mm_interconnect_1_hps_0_f2h_axi_slave_awvalid), //                   .awvalid
		.f2h_AWREADY                   (mm_interconnect_1_hps_0_f2h_axi_slave_awready), //                   .awready
		.f2h_AWUSER                    (mm_interconnect_1_hps_0_f2h_axi_slave_awuser),  //                   .awuser
		.f2h_WID                       (mm_interconnect_1_hps_0_f2h_axi_slave_wid),     //                   .wid
		.f2h_WDATA                     (mm_interconnect_1_hps_0_f2h_axi_slave_wdata),   //                   .wdata
		.f2h_WSTRB                     (mm_interconnect_1_hps_0_f2h_axi_slave_wstrb),   //                   .wstrb
		.f2h_WLAST                     (mm_interconnect_1_hps_0_f2h_axi_slave_wlast),   //                   .wlast
		.f2h_WVALID                    (mm_interconnect_1_hps_0_f2h_axi_slave_wvalid),  //                   .wvalid
		.f2h_WREADY                    (mm_interconnect_1_hps_0_f2h_axi_slave_wready),  //                   .wready
		.f2h_BID                       (mm_interconnect_1_hps_0_f2h_axi_slave_bid),     //                   .bid
		.f2h_BRESP                     (mm_interconnect_1_hps_0_f2h_axi_slave_bresp),   //                   .bresp
		.f2h_BVALID                    (mm_interconnect_1_hps_0_f2h_axi_slave_bvalid),  //                   .bvalid
		.f2h_BREADY                    (mm_interconnect_1_hps_0_f2h_axi_slave_bready),  //                   .bready
		.f2h_ARID                      (mm_interconnect_1_hps_0_f2h_axi_slave_arid),    //                   .arid
		.f2h_ARADDR                    (mm_interconnect_1_hps_0_f2h_axi_slave_araddr),  //                   .araddr
		.f2h_ARLEN                     (mm_interconnect_1_hps_0_f2h_axi_slave_arlen),   //                   .arlen
		.f2h_ARSIZE                    (mm_interconnect_1_hps_0_f2h_axi_slave_arsize),  //                   .arsize
		.f2h_ARBURST                   (mm_interconnect_1_hps_0_f2h_axi_slave_arburst), //                   .arburst
		.f2h_ARLOCK                    (mm_interconnect_1_hps_0_f2h_axi_slave_arlock),  //                   .arlock
		.f2h_ARCACHE                   (mm_interconnect_1_hps_0_f2h_axi_slave_arcache), //                   .arcache
		.f2h_ARPROT                    (mm_interconnect_1_hps_0_f2h_axi_slave_arprot),  //                   .arprot
		.f2h_ARVALID                   (mm_interconnect_1_hps_0_f2h_axi_slave_arvalid), //                   .arvalid
		.f2h_ARREADY                   (mm_interconnect_1_hps_0_f2h_axi_slave_arready), //                   .arready
		.f2h_ARUSER                    (mm_interconnect_1_hps_0_f2h_axi_slave_aruser),  //                   .aruser
		.f2h_RID                       (mm_interconnect_1_hps_0_f2h_axi_slave_rid),     //                   .rid
		.f2h_RDATA                     (mm_interconnect_1_hps_0_f2h_axi_slave_rdata),   //                   .rdata
		.f2h_RRESP                     (mm_interconnect_1_hps_0_f2h_axi_slave_rresp),   //                   .rresp
		.f2h_RLAST                     (mm_interconnect_1_hps_0_f2h_axi_slave_rlast),   //                   .rlast
		.f2h_RVALID                    (mm_interconnect_1_hps_0_f2h_axi_slave_rvalid),  //                   .rvalid
		.f2h_RREADY                    (mm_interconnect_1_hps_0_f2h_axi_slave_rready),  //                   .rready
		.h2f_lw_axi_clk                (clk_clk),                                       //   h2f_lw_axi_clock.clk
		.h2f_lw_AWID                   (hps_0_h2f_lw_axi_master_awid),                  //  h2f_lw_axi_master.awid
		.h2f_lw_AWADDR                 (hps_0_h2f_lw_axi_master_awaddr),                //                   .awaddr
		.h2f_lw_AWLEN                  (hps_0_h2f_lw_axi_master_awlen),                 //                   .awlen
		.h2f_lw_AWSIZE                 (hps_0_h2f_lw_axi_master_awsize),                //                   .awsize
		.h2f_lw_AWBURST                (hps_0_h2f_lw_axi_master_awburst),               //                   .awburst
		.h2f_lw_AWLOCK                 (hps_0_h2f_lw_axi_master_awlock),                //                   .awlock
		.h2f_lw_AWCACHE                (hps_0_h2f_lw_axi_master_awcache),               //                   .awcache
		.h2f_lw_AWPROT                 (hps_0_h2f_lw_axi_master_awprot),                //                   .awprot
		.h2f_lw_AWVALID                (hps_0_h2f_lw_axi_master_awvalid),               //                   .awvalid
		.h2f_lw_AWREADY                (hps_0_h2f_lw_axi_master_awready),               //                   .awready
		.h2f_lw_WID                    (hps_0_h2f_lw_axi_master_wid),                   //                   .wid
		.h2f_lw_WDATA                  (hps_0_h2f_lw_axi_master_wdata),                 //                   .wdata
		.h2f_lw_WSTRB                  (hps_0_h2f_lw_axi_master_wstrb),                 //                   .wstrb
		.h2f_lw_WLAST                  (hps_0_h2f_lw_axi_master_wlast),                 //                   .wlast
		.h2f_lw_WVALID                 (hps_0_h2f_lw_axi_master_wvalid),                //                   .wvalid
		.h2f_lw_WREADY                 (hps_0_h2f_lw_axi_master_wready),                //                   .wready
		.h2f_lw_BID                    (hps_0_h2f_lw_axi_master_bid),                   //                   .bid
		.h2f_lw_BRESP                  (hps_0_h2f_lw_axi_master_bresp),                 //                   .bresp
		.h2f_lw_BVALID                 (hps_0_h2f_lw_axi_master_bvalid),                //                   .bvalid
		.h2f_lw_BREADY                 (hps_0_h2f_lw_axi_master_bready),                //                   .bready
		.h2f_lw_ARID                   (hps_0_h2f_lw_axi_master_arid),                  //                   .arid
		.h2f_lw_ARADDR                 (hps_0_h2f_lw_axi_master_araddr),                //                   .araddr
		.h2f_lw_ARLEN                  (hps_0_h2f_lw_axi_master_arlen),                 //                   .arlen
		.h2f_lw_ARSIZE                 (hps_0_h2f_lw_axi_master_arsize),                //                   .arsize
		.h2f_lw_ARBURST                (hps_0_h2f_lw_axi_master_arburst),               //                   .arburst
		.h2f_lw_ARLOCK                 (hps_0_h2f_lw_axi_master_arlock),                //                   .arlock
		.h2f_lw_ARCACHE                (hps_0_h2f_lw_axi_master_arcache),               //                   .arcache
		.h2f_lw_ARPROT                 (hps_0_h2f_lw_axi_master_arprot),                //                   .arprot
		.h2f_lw_ARVALID                (hps_0_h2f_lw_axi_master_arvalid),               //                   .arvalid
		.h2f_lw_ARREADY                (hps_0_h2f_lw_axi_master_arready),               //                   .arready
		.h2f_lw_RID                    (hps_0_h2f_lw_axi_master_rid),                   //                   .rid
		.h2f_lw_RDATA                  (hps_0_h2f_lw_axi_master_rdata),                 //                   .rdata
		.h2f_lw_RRESP                  (hps_0_h2f_lw_axi_master_rresp),                 //                   .rresp
		.h2f_lw_RLAST                  (hps_0_h2f_lw_axi_master_rlast),                 //                   .rlast
		.h2f_lw_RVALID                 (hps_0_h2f_lw_axi_master_rvalid),                //                   .rvalid
		.h2f_lw_RREADY                 (hps_0_h2f_lw_axi_master_rready),                //                   .rready
		.f2h_irq_p0                    (hps_0_f2h_irq0_irq),                            //           f2h_irq0.irq
		.f2h_irq_p1                    (hps_0_f2h_irq1_irq)                             //           f2h_irq1.irq
	);

	i2c_opencores i2c_opencores_camera (
		.wb_clk_i   (clk_clk),                                                           //            clock.clk
		.wb_rst_i   (rst_controller_001_reset_out_reset),                                //      clock_reset.reset
		.scl_pad_io (i2c_opencores_camera_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_camera_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  ()                                                                   // interrupt_sender.irq
	);

	i2c_opencores i2c_opencores_mipi (
		.wb_clk_i   (clk_clk),                                                         //            clock.clk
		.wb_rst_i   (rst_controller_001_reset_out_reset),                              //      clock_reset.reset
		.scl_pad_io (i2c_opencores_mipi_export_scl_pad_io),                            //           export.export
		.sda_pad_io (i2c_opencores_mipi_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  ()                                                                 // interrupt_sender.irq
	);

	intr_capturer #(
		.NUM_INTR (32)
	) intr_capturer_0 (
		.clk          (clk_clk),                                                   //              clock.clk
		.rst_n        (~rst_controller_001_reset_out_reset),                       //         reset_sink.reset_n
		.addr         (mm_interconnect_3_intr_capturer_0_avalon_slave_0_address),  //     avalon_slave_0.address
		.read         (mm_interconnect_3_intr_capturer_0_avalon_slave_0_read),     //                   .read
		.rddata       (mm_interconnect_3_intr_capturer_0_avalon_slave_0_readdata), //                   .readdata
		.interrupt_in (intr_capturer_0_interrupt_receiver_irq)                     // interrupt_receiver.irq
	);

	soc_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_3_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_3_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_3_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_3_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_3_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_3_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_3_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	soc_system_key key (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_3_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)             //                 irq.irq
	);

	soc_system_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_3_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	soc_system_master_non_sec #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_non_sec (
		.clk_clk              (clk_clk),                             //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                      //    clk_reset.reset
		.master_address       (master_non_sec_master_address),       //       master.address
		.master_readdata      (master_non_sec_master_readdata),      //             .readdata
		.master_read          (master_non_sec_master_read),          //             .read
		.master_write         (master_non_sec_master_write),         //             .write
		.master_writedata     (master_non_sec_master_writedata),     //             .writedata
		.master_waitrequest   (master_non_sec_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_non_sec_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_non_sec_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                     // master_reset.reset
	);

	soc_system_master_non_sec #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_secure (
		.clk_clk              (clk_clk),                            //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                     //    clk_reset.reset
		.master_address       (master_secure_master_address),       //       master.address
		.master_readdata      (master_secure_master_readdata),      //             .readdata
		.master_read          (master_secure_master_read),          //             .read
		.master_write         (master_secure_master_write),         //             .write
		.master_writedata     (master_secure_master_writedata),     //             .writedata
		.master_waitrequest   (master_secure_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_secure_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_secure_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                    // master_reset.reset
	);

	soc_system_mipi_pwdn_n mipi_pwdn_n (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_3_mipi_pwdn_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_mipi_pwdn_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_mipi_pwdn_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_mipi_pwdn_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_mipi_pwdn_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_pwdn_n_external_connection_export)       // external_connection.export
	);

	soc_system_mipi_pwdn_n mipi_reset_n (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_3_mipi_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_mipi_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_mipi_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_mipi_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_mipi_reset_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_reset_n_external_connection_export)       // external_connection.export
	);

	soc_system_onchip_memory onchip_memory (
		.address     (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_2_onchip_memory_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_2_onchip_memory_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_2_onchip_memory_s2_clken),      //       .clken
		.write2      (mm_interconnect_2_onchip_memory_s2_write),      //       .write
		.readdata2   (mm_interconnect_2_onchip_memory_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_2_onchip_memory_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_2_onchip_memory_s2_byteenable), //       .byteenable
		.clk         (pll_0_outclk0_clk),                             //   clk1.clk
		.reset       (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	soc_system_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.outclk_1 (clk_sdram_clk),     // outclk1.clk
		.outclk_2 (d8m_xclkin_clk),    // outclk2.clk
		.outclk_3 (clk_vga_clk),       // outclk3.clk
		.locked   ()                   // (terminated)
	);

	soc_system_sdram sdram (
		.clk            (pll_0_outclk0_clk),                        //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_2_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_2_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_2_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_2_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_2_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_2_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_2_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_2_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_2_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	soc_system_st_adapter_0 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) st_adapter_0 (
		.in_clk_0_clk        (pll_0_outclk0_clk),                 // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),    // in_rst_0.reset
		.in_0_data           (alt_vip_cpr_2_dout1_data),          //     in_0.data
		.in_0_valid          (alt_vip_cpr_2_dout1_valid),         //         .valid
		.in_0_ready          (alt_vip_cpr_2_dout1_ready),         //         .ready
		.in_0_startofpacket  (alt_vip_cpr_2_dout1_startofpacket), //         .startofpacket
		.in_0_endofpacket    (alt_vip_cpr_2_dout1_endofpacket),   //         .endofpacket
		.out_0_data          (st_adapter_0_out_0_data),           //    out_0.data
		.out_0_valid         (st_adapter_0_out_0_valid),          //         .valid
		.out_0_ready         (st_adapter_0_out_0_ready),          //         .ready
		.out_0_startofpacket (st_adapter_0_out_0_startofpacket),  //         .startofpacket
		.out_0_endofpacket   (st_adapter_0_out_0_endofpacket)     //         .endofpacket
	);

	soc_system_sw sw (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_3_sw_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_3_sw_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_3_sw_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_3_sw_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_3_sw_s1_readdata),    //                    .readdata
		.in_port    (sw_external_connection_export),       // external_connection.export
		.irq        (irq_mapper_receiver2_irq)             //                 irq.irq
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_3_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_3_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_video_csc_0 video_csc_0 (
		.clk                      (pll_0_outclk0_clk),                           //               clk.clk
		.reset                    (rst_controller_reset_out_reset),              //             reset.reset
		.stream_in_startofpacket  (st_adapter_0_out_0_startofpacket),            //   avalon_csc_sink.startofpacket
		.stream_in_endofpacket    (st_adapter_0_out_0_endofpacket),              //                  .endofpacket
		.stream_in_valid          (st_adapter_0_out_0_valid),                    //                  .valid
		.stream_in_ready          (st_adapter_0_out_0_ready),                    //                  .ready
		.stream_in_data           (st_adapter_0_out_0_data),                     //                  .data
		.stream_out_ready         (video_csc_0_avalon_csc_source_ready),         // avalon_csc_source.ready
		.stream_out_startofpacket (video_csc_0_avalon_csc_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (video_csc_0_avalon_csc_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (video_csc_0_avalon_csc_source_valid),         //                  .valid
		.stream_out_data          (video_csc_0_avalon_csc_source_data)           //                  .data
	);

	soc_system_video_dma_controller_0 video_dma_controller_0 (
		.clk                  (pll_0_outclk0_clk),                                                            //                      clk.clk
		.reset                (rst_controller_reset_out_reset),                                               //                    reset.reset
		.stream_data          (video_csc_0_avalon_csc_source_data),                                           //          avalon_dma_sink.data
		.stream_startofpacket (video_csc_0_avalon_csc_source_startofpacket),                                  //                         .startofpacket
		.stream_endofpacket   (video_csc_0_avalon_csc_source_endofpacket),                                    //                         .endofpacket
		.stream_valid         (video_csc_0_avalon_csc_source_valid),                                          //                         .valid
		.stream_ready         (video_csc_0_avalon_csc_source_ready),                                          //                         .ready
		.slave_address        (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_readdata),   //                         .readdata
		.master_address       (video_dma_controller_0_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (video_dma_controller_0_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_write         (video_dma_controller_0_avalon_dma_master_write),                               //                         .write
		.master_writedata     (video_dma_controller_0_avalon_dma_master_writedata)                            //                         .writedata
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                                        (pll_0_outclk0_clk),                                    //                                      pll_0_outclk0.clk
		.video_dma_controller_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // video_dma_controller_0_reset_reset_bridge_in_reset.reset
		.video_dma_controller_0_avalon_dma_master_address         (video_dma_controller_0_avalon_dma_master_address),     //           video_dma_controller_0_avalon_dma_master.address
		.video_dma_controller_0_avalon_dma_master_waitrequest     (video_dma_controller_0_avalon_dma_master_waitrequest), //                                                   .waitrequest
		.video_dma_controller_0_avalon_dma_master_write           (video_dma_controller_0_avalon_dma_master_write),       //                                                   .write
		.video_dma_controller_0_avalon_dma_master_writedata       (video_dma_controller_0_avalon_dma_master_writedata),   //                                                   .writedata
		.onchip_memory_s1_address                                 (mm_interconnect_0_onchip_memory_s1_address),           //                                   onchip_memory_s1.address
		.onchip_memory_s1_write                                   (mm_interconnect_0_onchip_memory_s1_write),             //                                                   .write
		.onchip_memory_s1_readdata                                (mm_interconnect_0_onchip_memory_s1_readdata),          //                                                   .readdata
		.onchip_memory_s1_writedata                               (mm_interconnect_0_onchip_memory_s1_writedata),         //                                                   .writedata
		.onchip_memory_s1_byteenable                              (mm_interconnect_0_onchip_memory_s1_byteenable),        //                                                   .byteenable
		.onchip_memory_s1_chipselect                              (mm_interconnect_0_onchip_memory_s1_chipselect),        //                                                   .chipselect
		.onchip_memory_s1_clken                                   (mm_interconnect_0_onchip_memory_s1_clken)              //                                                   .clken
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_f2h_axi_slave_awid                                          (mm_interconnect_1_hps_0_f2h_axi_slave_awid),    //                                         hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                        (mm_interconnect_1_hps_0_f2h_axi_slave_awaddr),  //                                                            .awaddr
		.hps_0_f2h_axi_slave_awlen                                         (mm_interconnect_1_hps_0_f2h_axi_slave_awlen),   //                                                            .awlen
		.hps_0_f2h_axi_slave_awsize                                        (mm_interconnect_1_hps_0_f2h_axi_slave_awsize),  //                                                            .awsize
		.hps_0_f2h_axi_slave_awburst                                       (mm_interconnect_1_hps_0_f2h_axi_slave_awburst), //                                                            .awburst
		.hps_0_f2h_axi_slave_awlock                                        (mm_interconnect_1_hps_0_f2h_axi_slave_awlock),  //                                                            .awlock
		.hps_0_f2h_axi_slave_awcache                                       (mm_interconnect_1_hps_0_f2h_axi_slave_awcache), //                                                            .awcache
		.hps_0_f2h_axi_slave_awprot                                        (mm_interconnect_1_hps_0_f2h_axi_slave_awprot),  //                                                            .awprot
		.hps_0_f2h_axi_slave_awuser                                        (mm_interconnect_1_hps_0_f2h_axi_slave_awuser),  //                                                            .awuser
		.hps_0_f2h_axi_slave_awvalid                                       (mm_interconnect_1_hps_0_f2h_axi_slave_awvalid), //                                                            .awvalid
		.hps_0_f2h_axi_slave_awready                                       (mm_interconnect_1_hps_0_f2h_axi_slave_awready), //                                                            .awready
		.hps_0_f2h_axi_slave_wid                                           (mm_interconnect_1_hps_0_f2h_axi_slave_wid),     //                                                            .wid
		.hps_0_f2h_axi_slave_wdata                                         (mm_interconnect_1_hps_0_f2h_axi_slave_wdata),   //                                                            .wdata
		.hps_0_f2h_axi_slave_wstrb                                         (mm_interconnect_1_hps_0_f2h_axi_slave_wstrb),   //                                                            .wstrb
		.hps_0_f2h_axi_slave_wlast                                         (mm_interconnect_1_hps_0_f2h_axi_slave_wlast),   //                                                            .wlast
		.hps_0_f2h_axi_slave_wvalid                                        (mm_interconnect_1_hps_0_f2h_axi_slave_wvalid),  //                                                            .wvalid
		.hps_0_f2h_axi_slave_wready                                        (mm_interconnect_1_hps_0_f2h_axi_slave_wready),  //                                                            .wready
		.hps_0_f2h_axi_slave_bid                                           (mm_interconnect_1_hps_0_f2h_axi_slave_bid),     //                                                            .bid
		.hps_0_f2h_axi_slave_bresp                                         (mm_interconnect_1_hps_0_f2h_axi_slave_bresp),   //                                                            .bresp
		.hps_0_f2h_axi_slave_bvalid                                        (mm_interconnect_1_hps_0_f2h_axi_slave_bvalid),  //                                                            .bvalid
		.hps_0_f2h_axi_slave_bready                                        (mm_interconnect_1_hps_0_f2h_axi_slave_bready),  //                                                            .bready
		.hps_0_f2h_axi_slave_arid                                          (mm_interconnect_1_hps_0_f2h_axi_slave_arid),    //                                                            .arid
		.hps_0_f2h_axi_slave_araddr                                        (mm_interconnect_1_hps_0_f2h_axi_slave_araddr),  //                                                            .araddr
		.hps_0_f2h_axi_slave_arlen                                         (mm_interconnect_1_hps_0_f2h_axi_slave_arlen),   //                                                            .arlen
		.hps_0_f2h_axi_slave_arsize                                        (mm_interconnect_1_hps_0_f2h_axi_slave_arsize),  //                                                            .arsize
		.hps_0_f2h_axi_slave_arburst                                       (mm_interconnect_1_hps_0_f2h_axi_slave_arburst), //                                                            .arburst
		.hps_0_f2h_axi_slave_arlock                                        (mm_interconnect_1_hps_0_f2h_axi_slave_arlock),  //                                                            .arlock
		.hps_0_f2h_axi_slave_arcache                                       (mm_interconnect_1_hps_0_f2h_axi_slave_arcache), //                                                            .arcache
		.hps_0_f2h_axi_slave_arprot                                        (mm_interconnect_1_hps_0_f2h_axi_slave_arprot),  //                                                            .arprot
		.hps_0_f2h_axi_slave_aruser                                        (mm_interconnect_1_hps_0_f2h_axi_slave_aruser),  //                                                            .aruser
		.hps_0_f2h_axi_slave_arvalid                                       (mm_interconnect_1_hps_0_f2h_axi_slave_arvalid), //                                                            .arvalid
		.hps_0_f2h_axi_slave_arready                                       (mm_interconnect_1_hps_0_f2h_axi_slave_arready), //                                                            .arready
		.hps_0_f2h_axi_slave_rid                                           (mm_interconnect_1_hps_0_f2h_axi_slave_rid),     //                                                            .rid
		.hps_0_f2h_axi_slave_rdata                                         (mm_interconnect_1_hps_0_f2h_axi_slave_rdata),   //                                                            .rdata
		.hps_0_f2h_axi_slave_rresp                                         (mm_interconnect_1_hps_0_f2h_axi_slave_rresp),   //                                                            .rresp
		.hps_0_f2h_axi_slave_rlast                                         (mm_interconnect_1_hps_0_f2h_axi_slave_rlast),   //                                                            .rlast
		.hps_0_f2h_axi_slave_rvalid                                        (mm_interconnect_1_hps_0_f2h_axi_slave_rvalid),  //                                                            .rvalid
		.hps_0_f2h_axi_slave_rready                                        (mm_interconnect_1_hps_0_f2h_axi_slave_rready),  //                                                            .rready
		.clk_0_clk_clk                                                     (clk_clk),                                       //                                                   clk_0_clk.clk
		.pll_0_outclk0_clk                                                 (pll_0_outclk0_clk),                             //                                               pll_0_outclk0.clk
		.alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                //    alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset.reset
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset  (rst_controller_002_reset_out_reset),            //  hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.master_secure_clk_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),            //               master_secure_clk_reset_reset_bridge_in_reset.reset
		.master_secure_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),            // master_secure_master_translator_reset_reset_bridge_in_reset.reset
		.alt_vip_vfr_vga_avalon_master_address                             (alt_vip_vfr_vga_avalon_master_address),         //                               alt_vip_vfr_vga_avalon_master.address
		.alt_vip_vfr_vga_avalon_master_waitrequest                         (alt_vip_vfr_vga_avalon_master_waitrequest),     //                                                            .waitrequest
		.alt_vip_vfr_vga_avalon_master_burstcount                          (alt_vip_vfr_vga_avalon_master_burstcount),      //                                                            .burstcount
		.alt_vip_vfr_vga_avalon_master_read                                (alt_vip_vfr_vga_avalon_master_read),            //                                                            .read
		.alt_vip_vfr_vga_avalon_master_readdata                            (alt_vip_vfr_vga_avalon_master_readdata),        //                                                            .readdata
		.alt_vip_vfr_vga_avalon_master_readdatavalid                       (alt_vip_vfr_vga_avalon_master_readdatavalid),   //                                                            .readdatavalid
		.master_secure_master_address                                      (master_secure_master_address),                  //                                        master_secure_master.address
		.master_secure_master_waitrequest                                  (master_secure_master_waitrequest),              //                                                            .waitrequest
		.master_secure_master_byteenable                                   (master_secure_master_byteenable),               //                                                            .byteenable
		.master_secure_master_read                                         (master_secure_master_read),                     //                                                            .read
		.master_secure_master_readdata                                     (master_secure_master_readdata),                 //                                                            .readdata
		.master_secure_master_readdatavalid                                (master_secure_master_readdatavalid),            //                                                            .readdatavalid
		.master_secure_master_write                                        (master_secure_master_write),                    //                                                            .write
		.master_secure_master_writedata                                    (master_secure_master_writedata)                 //                                                            .writedata
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                     //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                   //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                    //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                   //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                  //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                   //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                  //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                   //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                  //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                  //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                      //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                    //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                    //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                    //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                   //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                   //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                      //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                    //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                   //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                   //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                     //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                   //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                    //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                   //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                  //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                   //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                  //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                   //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                  //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                  //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                      //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                    //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                    //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                    //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                   //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                   //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                       //                                                  clk_0_clk.clk
		.pll_0_outclk0_clk                                                (pll_0_outclk0_clk),                             //                                              pll_0_outclk0.clk
		.alt_vip_vfb_0_reset_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                //                  alt_vip_vfb_0_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),            // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.alt_vip_vfb_0_read_master_address                                (alt_vip_vfb_0_read_master_address),             //                                  alt_vip_vfb_0_read_master.address
		.alt_vip_vfb_0_read_master_waitrequest                            (alt_vip_vfb_0_read_master_waitrequest),         //                                                           .waitrequest
		.alt_vip_vfb_0_read_master_burstcount                             (alt_vip_vfb_0_read_master_burstcount),          //                                                           .burstcount
		.alt_vip_vfb_0_read_master_read                                   (alt_vip_vfb_0_read_master_read),                //                                                           .read
		.alt_vip_vfb_0_read_master_readdata                               (alt_vip_vfb_0_read_master_readdata),            //                                                           .readdata
		.alt_vip_vfb_0_read_master_readdatavalid                          (alt_vip_vfb_0_read_master_readdatavalid),       //                                                           .readdatavalid
		.alt_vip_vfb_0_write_master_address                               (alt_vip_vfb_0_write_master_address),            //                                 alt_vip_vfb_0_write_master.address
		.alt_vip_vfb_0_write_master_waitrequest                           (alt_vip_vfb_0_write_master_waitrequest),        //                                                           .waitrequest
		.alt_vip_vfb_0_write_master_burstcount                            (alt_vip_vfb_0_write_master_burstcount),         //                                                           .burstcount
		.alt_vip_vfb_0_write_master_write                                 (alt_vip_vfb_0_write_master_write),              //                                                           .write
		.alt_vip_vfb_0_write_master_writedata                             (alt_vip_vfb_0_write_master_writedata),          //                                                           .writedata
		.onchip_memory_s2_address                                         (mm_interconnect_2_onchip_memory_s2_address),    //                                           onchip_memory_s2.address
		.onchip_memory_s2_write                                           (mm_interconnect_2_onchip_memory_s2_write),      //                                                           .write
		.onchip_memory_s2_readdata                                        (mm_interconnect_2_onchip_memory_s2_readdata),   //                                                           .readdata
		.onchip_memory_s2_writedata                                       (mm_interconnect_2_onchip_memory_s2_writedata),  //                                                           .writedata
		.onchip_memory_s2_byteenable                                      (mm_interconnect_2_onchip_memory_s2_byteenable), //                                                           .byteenable
		.onchip_memory_s2_chipselect                                      (mm_interconnect_2_onchip_memory_s2_chipselect), //                                                           .chipselect
		.onchip_memory_s2_clken                                           (mm_interconnect_2_onchip_memory_s2_clken),      //                                                           .clken
		.sdram_s1_address                                                 (mm_interconnect_2_sdram_s1_address),            //                                                   sdram_s1.address
		.sdram_s1_write                                                   (mm_interconnect_2_sdram_s1_write),              //                                                           .write
		.sdram_s1_read                                                    (mm_interconnect_2_sdram_s1_read),               //                                                           .read
		.sdram_s1_readdata                                                (mm_interconnect_2_sdram_s1_readdata),           //                                                           .readdata
		.sdram_s1_writedata                                               (mm_interconnect_2_sdram_s1_writedata),          //                                                           .writedata
		.sdram_s1_byteenable                                              (mm_interconnect_2_sdram_s1_byteenable),         //                                                           .byteenable
		.sdram_s1_readdatavalid                                           (mm_interconnect_2_sdram_s1_readdatavalid),      //                                                           .readdatavalid
		.sdram_s1_waitrequest                                             (mm_interconnect_2_sdram_s1_waitrequest),        //                                                           .waitrequest
		.sdram_s1_chipselect                                              (mm_interconnect_2_sdram_s1_chipselect)          //                                                           .chipselect
	);

	soc_system_mm_interconnect_3 mm_interconnect_3 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                                 //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                                               //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                                                //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                                               //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                                              //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                                               //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                                              //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                                               //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                                              //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                                              //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                                  //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                                                //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                                                //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                                                //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                                               //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                                               //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                                  //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                                                //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                                               //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                                               //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                                 //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                                               //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                                                //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                                               //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                                              //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                                               //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                                              //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                                               //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                                              //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                                              //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                                  //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                                                //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                                                //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                                                //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                                               //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                                               //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                                      //                                                     clk_0_clk.clk
		.pll_0_outclk0_clk                                                   (pll_0_outclk0_clk),                                                            //                                                 pll_0_outclk0.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                           // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset                         (rst_controller_001_reset_out_reset),                                           //                         jtag_uart_reset_reset_bridge_in_reset.reset
		.master_non_sec_clk_reset_reset_bridge_in_reset_reset                (rst_controller_001_reset_out_reset),                                           //                master_non_sec_clk_reset_reset_bridge_in_reset.reset
		.video_dma_controller_0_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                                               //            video_dma_controller_0_reset_reset_bridge_in_reset.reset
		.master_non_sec_master_address                                       (master_non_sec_master_address),                                                //                                         master_non_sec_master.address
		.master_non_sec_master_waitrequest                                   (master_non_sec_master_waitrequest),                                            //                                                              .waitrequest
		.master_non_sec_master_byteenable                                    (master_non_sec_master_byteenable),                                             //                                                              .byteenable
		.master_non_sec_master_read                                          (master_non_sec_master_read),                                                   //                                                              .read
		.master_non_sec_master_readdata                                      (master_non_sec_master_readdata),                                               //                                                              .readdata
		.master_non_sec_master_readdatavalid                                 (master_non_sec_master_readdatavalid),                                          //                                                              .readdatavalid
		.master_non_sec_master_write                                         (master_non_sec_master_write),                                                  //                                                              .write
		.master_non_sec_master_writedata                                     (master_non_sec_master_writedata),                                              //                                                              .writedata
		.alt_vip_cl_clp_1_control_address                                    (mm_interconnect_3_alt_vip_cl_clp_1_control_address),                           //                                      alt_vip_cl_clp_1_control.address
		.alt_vip_cl_clp_1_control_write                                      (mm_interconnect_3_alt_vip_cl_clp_1_control_write),                             //                                                              .write
		.alt_vip_cl_clp_1_control_read                                       (mm_interconnect_3_alt_vip_cl_clp_1_control_read),                              //                                                              .read
		.alt_vip_cl_clp_1_control_readdata                                   (mm_interconnect_3_alt_vip_cl_clp_1_control_readdata),                          //                                                              .readdata
		.alt_vip_cl_clp_1_control_writedata                                  (mm_interconnect_3_alt_vip_cl_clp_1_control_writedata),                         //                                                              .writedata
		.alt_vip_cl_clp_1_control_byteenable                                 (mm_interconnect_3_alt_vip_cl_clp_1_control_byteenable),                        //                                                              .byteenable
		.alt_vip_cl_clp_1_control_readdatavalid                              (mm_interconnect_3_alt_vip_cl_clp_1_control_readdatavalid),                     //                                                              .readdatavalid
		.alt_vip_cl_clp_1_control_waitrequest                                (mm_interconnect_3_alt_vip_cl_clp_1_control_waitrequest),                       //                                                              .waitrequest
		.alt_vip_mix_0_control_address                                       (mm_interconnect_3_alt_vip_mix_0_control_address),                              //                                         alt_vip_mix_0_control.address
		.alt_vip_mix_0_control_write                                         (mm_interconnect_3_alt_vip_mix_0_control_write),                                //                                                              .write
		.alt_vip_mix_0_control_readdata                                      (mm_interconnect_3_alt_vip_mix_0_control_readdata),                             //                                                              .readdata
		.alt_vip_mix_0_control_writedata                                     (mm_interconnect_3_alt_vip_mix_0_control_writedata),                            //                                                              .writedata
		.alt_vip_mix_0_control_chipselect                                    (mm_interconnect_3_alt_vip_mix_0_control_chipselect),                           //                                                              .chipselect
		.alt_vip_vfr_vga_avalon_slave_address                                (mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_address),                       //                                  alt_vip_vfr_vga_avalon_slave.address
		.alt_vip_vfr_vga_avalon_slave_write                                  (mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_write),                         //                                                              .write
		.alt_vip_vfr_vga_avalon_slave_read                                   (mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_read),                          //                                                              .read
		.alt_vip_vfr_vga_avalon_slave_readdata                               (mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_readdata),                      //                                                              .readdata
		.alt_vip_vfr_vga_avalon_slave_writedata                              (mm_interconnect_3_alt_vip_vfr_vga_avalon_slave_writedata),                     //                                                              .writedata
		.i2c_opencores_camera_avalon_slave_0_address                         (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_address),                //                           i2c_opencores_camera_avalon_slave_0.address
		.i2c_opencores_camera_avalon_slave_0_write                           (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_write),                  //                                                              .write
		.i2c_opencores_camera_avalon_slave_0_readdata                        (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_readdata),               //                                                              .readdata
		.i2c_opencores_camera_avalon_slave_0_writedata                       (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_writedata),              //                                                              .writedata
		.i2c_opencores_camera_avalon_slave_0_waitrequest                     (~mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_waitrequest),           //                                                              .waitrequest
		.i2c_opencores_camera_avalon_slave_0_chipselect                      (mm_interconnect_3_i2c_opencores_camera_avalon_slave_0_chipselect),             //                                                              .chipselect
		.i2c_opencores_mipi_avalon_slave_0_address                           (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_address),                  //                             i2c_opencores_mipi_avalon_slave_0.address
		.i2c_opencores_mipi_avalon_slave_0_write                             (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_write),                    //                                                              .write
		.i2c_opencores_mipi_avalon_slave_0_readdata                          (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_readdata),                 //                                                              .readdata
		.i2c_opencores_mipi_avalon_slave_0_writedata                         (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_writedata),                //                                                              .writedata
		.i2c_opencores_mipi_avalon_slave_0_waitrequest                       (~mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_waitrequest),             //                                                              .waitrequest
		.i2c_opencores_mipi_avalon_slave_0_chipselect                        (mm_interconnect_3_i2c_opencores_mipi_avalon_slave_0_chipselect),               //                                                              .chipselect
		.intr_capturer_0_avalon_slave_0_address                              (mm_interconnect_3_intr_capturer_0_avalon_slave_0_address),                     //                                intr_capturer_0_avalon_slave_0.address
		.intr_capturer_0_avalon_slave_0_read                                 (mm_interconnect_3_intr_capturer_0_avalon_slave_0_read),                        //                                                              .read
		.intr_capturer_0_avalon_slave_0_readdata                             (mm_interconnect_3_intr_capturer_0_avalon_slave_0_readdata),                    //                                                              .readdata
		.jtag_uart_avalon_jtag_slave_address                                 (mm_interconnect_3_jtag_uart_avalon_jtag_slave_address),                        //                                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                   (mm_interconnect_3_jtag_uart_avalon_jtag_slave_write),                          //                                                              .write
		.jtag_uart_avalon_jtag_slave_read                                    (mm_interconnect_3_jtag_uart_avalon_jtag_slave_read),                           //                                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                                (mm_interconnect_3_jtag_uart_avalon_jtag_slave_readdata),                       //                                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata                               (mm_interconnect_3_jtag_uart_avalon_jtag_slave_writedata),                      //                                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                             (mm_interconnect_3_jtag_uart_avalon_jtag_slave_waitrequest),                    //                                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                              (mm_interconnect_3_jtag_uart_avalon_jtag_slave_chipselect),                     //                                                              .chipselect
		.key_s1_address                                                      (mm_interconnect_3_key_s1_address),                                             //                                                        key_s1.address
		.key_s1_write                                                        (mm_interconnect_3_key_s1_write),                                               //                                                              .write
		.key_s1_readdata                                                     (mm_interconnect_3_key_s1_readdata),                                            //                                                              .readdata
		.key_s1_writedata                                                    (mm_interconnect_3_key_s1_writedata),                                           //                                                              .writedata
		.key_s1_chipselect                                                   (mm_interconnect_3_key_s1_chipselect),                                          //                                                              .chipselect
		.led_s1_address                                                      (mm_interconnect_3_led_s1_address),                                             //                                                        led_s1.address
		.led_s1_write                                                        (mm_interconnect_3_led_s1_write),                                               //                                                              .write
		.led_s1_readdata                                                     (mm_interconnect_3_led_s1_readdata),                                            //                                                              .readdata
		.led_s1_writedata                                                    (mm_interconnect_3_led_s1_writedata),                                           //                                                              .writedata
		.led_s1_chipselect                                                   (mm_interconnect_3_led_s1_chipselect),                                          //                                                              .chipselect
		.mipi_pwdn_n_s1_address                                              (mm_interconnect_3_mipi_pwdn_n_s1_address),                                     //                                                mipi_pwdn_n_s1.address
		.mipi_pwdn_n_s1_write                                                (mm_interconnect_3_mipi_pwdn_n_s1_write),                                       //                                                              .write
		.mipi_pwdn_n_s1_readdata                                             (mm_interconnect_3_mipi_pwdn_n_s1_readdata),                                    //                                                              .readdata
		.mipi_pwdn_n_s1_writedata                                            (mm_interconnect_3_mipi_pwdn_n_s1_writedata),                                   //                                                              .writedata
		.mipi_pwdn_n_s1_chipselect                                           (mm_interconnect_3_mipi_pwdn_n_s1_chipselect),                                  //                                                              .chipselect
		.mipi_reset_n_s1_address                                             (mm_interconnect_3_mipi_reset_n_s1_address),                                    //                                               mipi_reset_n_s1.address
		.mipi_reset_n_s1_write                                               (mm_interconnect_3_mipi_reset_n_s1_write),                                      //                                                              .write
		.mipi_reset_n_s1_readdata                                            (mm_interconnect_3_mipi_reset_n_s1_readdata),                                   //                                                              .readdata
		.mipi_reset_n_s1_writedata                                           (mm_interconnect_3_mipi_reset_n_s1_writedata),                                  //                                                              .writedata
		.mipi_reset_n_s1_chipselect                                          (mm_interconnect_3_mipi_reset_n_s1_chipselect),                                 //                                                              .chipselect
		.sw_s1_address                                                       (mm_interconnect_3_sw_s1_address),                                              //                                                         sw_s1.address
		.sw_s1_write                                                         (mm_interconnect_3_sw_s1_write),                                                //                                                              .write
		.sw_s1_readdata                                                      (mm_interconnect_3_sw_s1_readdata),                                             //                                                              .readdata
		.sw_s1_writedata                                                     (mm_interconnect_3_sw_s1_writedata),                                            //                                                              .writedata
		.sw_s1_chipselect                                                    (mm_interconnect_3_sw_s1_chipselect),                                           //                                                              .chipselect
		.sysid_qsys_control_slave_address                                    (mm_interconnect_3_sysid_qsys_control_slave_address),                           //                                      sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                                   (mm_interconnect_3_sysid_qsys_control_slave_readdata),                          //                                                              .readdata
		.video_dma_controller_0_avalon_dma_control_slave_address             (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_address),    //               video_dma_controller_0_avalon_dma_control_slave.address
		.video_dma_controller_0_avalon_dma_control_slave_write               (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_write),      //                                                              .write
		.video_dma_controller_0_avalon_dma_control_slave_read                (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_read),       //                                                              .read
		.video_dma_controller_0_avalon_dma_control_slave_readdata            (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_readdata),   //                                                              .readdata
		.video_dma_controller_0_avalon_dma_control_slave_writedata           (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_writedata),  //                                                              .writedata
		.video_dma_controller_0_avalon_dma_control_slave_byteenable          (mm_interconnect_3_video_dma_controller_0_avalon_dma_control_slave_byteenable)  //                                                              .byteenable
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_002 (
		.clk           (clk_clk),                                //       clk.clk
		.reset         (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),               // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),               // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),               // receiver2.irq
		.sender_irq    (intr_capturer_0_interrupt_receiver_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
