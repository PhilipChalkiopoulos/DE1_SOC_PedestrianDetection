��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�v<��m���X#�m�o*�����z5�22�8�G4�x�{[��IW��(X(_<A�&��աW�����T��)΅�A�P���)���0� #7><����r|ES[��~�D $:_R.`
Hաm[��B,�+�*	p�xX��$��e�����?���G��%Z��Ǟ�H� �a�C��|�� �P�'Ђ�����|o�]1��%���L��a�B�JN���9�k���yEoȈ Xͬ���j���*��y"F��Z�G�>�FR�+�j�*��u"�pސz�x�Z&<�x����.s��!
$SϸΉ��'�EX�l@L]�C��z(Ka/�C��Sv�-��%-b�}�`�x$c;�Jl�:��9�T�KCx�^�3��S��|�p�hp*��l]�KwBDU�ȣ����O� �k�Q"|�"p��v&xW��9�
؎Җ�����Q�y���p0���]���9g^�ڙ; �5�)��~Lo��9�����l]�k�m��Te-!�
\�K��#�,��͜[�頚���bڳk�Gj��=��Ɯ-�À�y�Xi���8�6{����5���/�M�ݛ���I�d�;�!�;���,��)#��> ��-���لM2����縏;����N�,�D*)��$��٧68��6A�bA�#�#� -�
C��!{q{�sz�c$Ň>}@{]���mO���YD��1Jl���\f��F+Z>k����7�6eɖ HK���2�.Z�5�xdދ���3N��_�a�SЗ��G� �+�^�d�v�s��gN�p�[�;�w���A���kȽ8��/S�׊ր�0��x^�(�DESy��T������D7��6Z�m0����
z�E�h"�+`s�V16}*���Q�Z>�{y�����
(S���jL%M��دݿVM��]WWA�vp��)�fb������w.+,��'�ǉwճ*xs*h
��� οj ���'��JWn�z�����'�q+����}WG�mT}2e���Sh�#5��B%&�0�@f�`�L
Spy��9JpH����\���G���o�����nޯt*�T�	j�D`2�z�9��L�A�^��Q�ɯW̃4A�gH��i���'��D�|��餦��3�������em��u�β�&�DPz�J�]5����W���6Xg�6�v.4���\����Kp�˥LkR��0���2�s]�EEWp����� pv��]���թb�V�Zա+�7��+$�PZ��!�k�rq|'�>Z������&��E0ﵨ6ǩj���*�&�ގ��Al�zh�v���ULc��)�)�QJ6z2V�S<�4t�7��6�o] И8=8
?e���ب��\i	�1�O�8xMz�R2�	3��|c�x�����w!R�d�[�,�|u�� �H]�ҹ���
��^�f��+;Hf7v���)s�%���ĵ����,�x�NA$�i� ���;�R�w�8Q�� ���F�����b��::���H*�j��G!]"@����e^ٗ1L������Ub�bdUU�¨���$�AL|/ѣ#��%�胨P�:`ve��Fz�ka���ePK���+��a�5|���<�|3�&��2�t'�z�`W="����`�]�G���L
���o'�7�Mu���NH���	=���Y�7sip,��~a�YI�O�*��F�������ܮ��(/2���n�ꠇyT�(E&D6��T�p&'|�ȑ��~"$s��� z�/o�c�����h��-F��F��l�A�����)�W���86�G��1,D0=/���C�OF@, �`�ީ,otTr��Q���C�7\�A�J�r5�ֿ��S��M�9`��k��\#�d��\3�:�m�"��G�(�G�ѵGY��{���zAA��~P Tδv��ZIxN�QM]#�
`����u�3
b������0v���s��"-@��)t�l�[[�
�@�F�:�c\w�O����� ��|����0a�b�F���������)�a��d�N�ꉻ'���~nЁ{��h&�:1�)p��)��(�u��=���"���)0�����ȴ�%�#�4���yf$jX#7ߴ�k�f��P�o��I��s�?<�(�����(}�Lu�)� ��j�i/u���:)$.b�[[�I���bw_v��z�)޽Q�hS��zsF���4!���|�*��|�e�s�%$T���V�<i{�֬\�����`�|*����$El	.1a�����H����uFj[F���p�X�RT�+���1�ee��@V��w�]u���#\��yD���|�E�~B�c�z$e
���8X#�v�l��}Y�
5Ճ�D0ɂi\\��
�siG��t�g��;�	h��I��*��_��1Ր��s��GE�$�1B�O��*����Z ������l;mvp�ӣ�?��� �{��Yk���YaV+�\��=��ݑ����\ͬ]�I�-�X,ϋ}�_Z6��O�)\�(���5,uPI��!g�f���/��e�����U}���P.�zūzS�l��u�{G9��!R�&Q#^�SP'(�����!f�
����nG\�>Z�G�:κ��W��.��c�q���w�a+�U��hI��uH�Z;~Sd0�;��!#��L��p ��͙�d�Ł�G���`_��˥�`)�G�j���*ǧi`d&��p=�wB��mS����w5;J���Q����K�<�v�.�m%\Jr1F�C~��9P�˴v��ǣ2A4d"�iV�)b��ӟ�稼���t����s���Qx��="�,M�t����o�p�6���l�H�?�MLF���*�v�q�b;��9���Ed�1�@CRU�����k����0��B],�	��q�0Wm���Md|B#��W��r��{�.�71M|=Ig��뻕�Vp-׮ Js2�SҼ
�&���N�K��XQ_c���gP�p��D����#4��9�D9=�Bị;��/��f$�7f�Y�K������t9\�9Ѥ�IA�Q��͓�Z�Z �^qC!ȇ������F$f;�4K;L��	2�AbI�����d���_�R���ZӠ�W�ñ�r�ݾ��jwD
��}�*��j��
�K�������!�;��?�cJ�7#���r�)-a;��x�Ւ��������೚24#gL���b��e~���ʿ��#l�w�9��_}�G]M ��� ����Ns�h���4BL��+�O����z�T����p�Ӂ�+�?�/9���Ќ�����X�~�+�ED��?�,v����&�߆�k��� �<�Tk�LdLr4V[D��Z5���uR2m5��v��.�>ŋH�מ� ����m�d�H�bM�#Eh{1�X�O�S���9@�����4�KL�)��'>��K����{�S5��B�q�~�B9�y,�}�AM�sl�,��%���3��y�X�6C���V$��h8�;��H�x6Wk�^���O|���;r+p ��8� i�@��i/��M�� �G�a��3�7��`��q$3�X�S�c�Y�p�7���Ecf��ϋͭ�س�y�2N�u��?a�X��2�+w�E�:^=L�.�C|�3q}=��Z���gX�{"� �ܖY��;�y�}|w�7w���(%ָ�:Xf�I�՗��u�8���?)�	;��y��#n�`T�|f�.�pmk�=F���A�4�%2�ţ|��>{��*�N����Ns�jUA���)��珧�(�#�q�݂>-�/�'
U��Q�*�?�L+��D�'�C[W�I�d�
 f"�$�T�+$��B�p��!�@%SX.���+}�DB4Α��r��j�Y�ֵW���dUO�Q��NT��1أ*牄Vq�u83��U��j�1i�� a�C༚��.r ����?>�۠j�����]�6�8ԧ�C/��r��j4y�׎_�h,M����6N�r��vfϖ^F���ە�pydƒ�E������{]!-e�ѡݸQ[�u�Z�'�H���[�A�����Ec_F^�����]<�T�;O%%�𥥳�}��+�<l��t���\��h�a�IGP�)o��wO$c�Ur^�Yk��ϭw�[�V��V_6�۰W��;y*�����9߹��S��I���=A ��cO5��k�Q�sɯWus�$*�����4o�'.�׉c�qɜ��N����d"xԭD�`�sY	�@�QY�4Tv�þ�zB��fGv����B��w� ^d 	�]���N�9�΢����2��#W��=�&=����"�Ǘٰ�-�Šj�c���͞[�r�q��5�����2<#Z�3Z�(e��~�R�q�Åw�q=c�go���/�6G�j�ny�#��A��Y3lv��2���Z�oC���C|�[��	���ճ��ƌq��{�H�Kk�+�s�y=�/�Up � p��QYo��:��q��,��S��L.�̩F��D�zఔ�*aXS h8?��wbR�e��E;�g��
��%G�<�+�|�)��K���p����sa7'j����=`��O�BV�@_2)dG�%!���^B���"g��[9��M]HH�0�l�=|W#�)���xm7=�������j�_2�䏦&M����W&���%抳�u����GEM�O>���2���L�>�]���O7!7�`��N��=$A��9���* ��f�敧�Ar#EdvϦ��Z����J=��tЅQ��Ec�@P���f,�$'h四Օ���t��8�_���="�h�;B�IE���Fm��Xr'��d3ҹHL�	�m���x�`cP��y��,_�D�q���?��K��k�0y�p���c�Mǘ*SO�B/�� `ɬ�a����y@����5a��+�vrd�a���>�N%�5;:�ɴ�E�T@�FI�����Xb��x��Y�5�����|(�g�cm�p,=qN';h�j�i�qa�ƶQ�x�U�œ$��Y���a�y�} Y:Ҧ�؟|R~4槄Dql� �N��R��~�1Wλ����Z�[A�D��(��6|���D���m�I,J�Z�J�p)�־��J����c'�3��
���
��TԲK�ە���6���*gU��]1fU�Ŵ���_���B�������Wn׃��ܫmR���l�M�����+!�y���`��1��G��%V������[��{T:E"_�!�F��6�� ��Ѐ��X��¾��Js�g��/��Z5�i�T���}�v
��.�����4Ǔ�n��[^Mm��=��>sp�;�f'MA���4L��N�#C����6�t%x�eS[�=>�M�d�w�ь���@S	#	vI,�9�>��M^R��a���x- @{��r���3C/��_|9I��>�V���[��֩�3 ��J����S�4��,�N�J�$)r|>^)�����y�j?���4��+�]�$C?Ɗ(��f^x��8�~ͦ!��[l~����s�v/t82�t!��iebf��3��`F#��#�ŀ�R*�^?�~��B\;*��Ƶz�ԬQQW��*C�ӷ���;t�49��¯�ˢ��6�.����.�N�<9����d��Tv۸r4ب��}�Y�6��d��Za����\#�'R�S�VF$�u]�*
}%\��~6��V���/��׻k����y4�x�I���[	XPR���z&����qw��~6iԱ�`���|I.�U����Sw���Mr�a�MP���މ��`�/�Xސ�F��ۏy�X��ʣ7���ڈh�?Mn%ؿ=^��i@�����`�u���|��K���ly��!�u�8�H~�gq��9	���Ϋ�|�-6">��F<�L���(��L��	���XX���u���N�2�Hi0
C�^��X�e�����]  NA�,�1�V�J���������	�0�e�jz:k�ZX��
� ����a�_��8�а��H�	��}.��f�_�C�x�-�;A1o�4a�It9�<�dmX�U!�QŠ �aMN�"��J��$��]+37��9��HE���`�����S��}�>*��2uσ~rj\�	J�t��v�`U_5{�������@��RE���Τw������E�8#��:аhf7P��F9�k7�Ю\	�>t�-	���ή��,�g|A�5��do�&ڒ�^��8G��ɕ0���F%l�L"�Ffp�:@�ŎBu�X!�[p2�`h��.��@c�	��Hrüt��Z1T�]���U�����g�XQ4yyU��B^A7	���J>Q��r.	��?�},����oYЅ'�y���*-���B�@�w��o �_~���"��e���qp����_��$ۦfjUh��Y�ag#ݞ���^�ք����bI�i~�J2�؜|���ׂ�,b��l���Wd$��> ��쬍�0�$�+���e��`� �a����;�{ϲ��,^p@mOh�|RA�`�U�"��B�/In����/�^���������S�8\�8V�x���r����T����4J�4����? @;�Dsb�,HQ�� �ߜ�7a;�~L��=p�q��E�,������QL�L���������q��8Mҫ�� ��Bh�{�1��?�O��t.�0�C�US|��:����Sp�J|ڼ
ꖍ3� �����R��*gmغ�
������0"��ub�o���j*#�@�D���<ee�3��X�=>`�ւG���<&d�N��6@M��(��<r���\s~ �y#�E��V�����Q9�����'fE��"˶�Z>��<�5O2��h�W�]�d�Y�<
��L�{�}��i�OϢ�i=����ׄ����t��Lʾ��s ������3���(
����e �K<����]�e0j2�I<����=O�^Pg���dP�m�����,������f��RZ����h~)6�t�tbK���l�nwr����p�&��ݒ:����#�p9a�L�-���iĲ@���	����������i,o�e�Z�5��pk�Z�ZG��̊z俎�
 g��ꊥgY�,fv�>���{ៀ,v��N��sb"�s)]3��X�J�m����Ա�u'�׹ڏ�Ke,�Q�k�i_uy�ТP��udwd�B�N%@03=��}�ux��'-,�� tR��휳������������v�c��@	�������u�R5}����V�	VX
d�@8����ne׌��$ԦO�.�L���9�1'3�٥�Q&�}KYZ,�r\�"�|Gq5Q	��9���ȼ�ZH�	D���|s"�|���dt��(MoHLeR��v�����5K�*y� �jY���f�Fw: C��jh��ĝ�E�d4w�*��3Ҏ�&y9ӊ����Ni\.�2?ݔ� ˫���?��*;靔�[���X!B���5�oqH��O�9x�E3�~�'��8	�_ڃ$�2+��w�C8���8�������P��
�Y�v��E��YG�3rs1c��:Ѩ���`���;�x y��&���<�H ��Ӹ^zݖ�4��q�*�`�8��H�j���qN��Dz�A4��˱Q�5߿�X��CT?�;�Y��7D�&	:[؛.(���,�{�3оt��!�K&��3;m8D�\�Iحb|_�v̼�? Rn7��Z�!��/��.!�{�\��F6���?G,_=j8�]��&S��x��^OM.��R'����G��@ ��`�wU��E7Ǉ"�[��;BN���� �� �����{8K��b�[��J0̐>yU�2]؝IBPy����3�NAp�ƹ<����۱���F؊t��IXk	�:�ƔpdY2��X唝}�"�ڪ��A��Id���_	8�,]���&�U�����6F�C��=�[�w7��؇������g��}���-�$`x���g���f�	ܗr9D�Lj�!?�C��T�ݎ�cP*��$��1X�ҧ�j��Jv�D�,�
��[�Ǡ��fg��`�B���`Vm�H��J���egm%f�է-��_s�����*�4�m�vky�'�
=�[�<�Τ�*�h������kki	(!2[(��FJ�b-1�]/���Y?�Ŧ��NSes $��ʞ���m�!K*��5م^��-�X��C�µԑ��Ĳ0�z�?�b�>zU�	}?z+T-A�A��҅h�p~�p3BGuU��y����21B]g��y��,���wۉH��&/���Cen�F!(J������%S�Ș���2q@E�*:�X�dl]�8(3�������Ӄy^&>}�-㰂c��k!z#�#�4)�S4�U|w<PA�IEE��:d�U&b��֊���2?��uR�o�KB)Q��%ލWm���Z�*m[=!u�Z���eZ��T\���nB ���֦F 	��g��F������OWK�W�v�D�R�����>7eYe;��t�Ꝓ��=��Zap�*!ʉU�~!q���	��ث�&�m~�qW6/v$��z�Pm,�!o-E�.��x�G 5c�Y����}5>���t֬C#�s���a��=K�\���D/Q1�V������$n�gs�g�ӹ#��TB����	�� .
V�Xn��C��1�z����ۊ��Ch��+����Jr�Ҽ$e�����������*O��%����r�ۓ���
T�A�"�&���l�m�#l�2�����^E���/��ʞ�T�TH���O���:���lnIˠ滬�3I����'A�*.>6���C!b%�fb�c�Q����&P$���_�k��?kC��怄�6&���|�Iw���8|]l�&N��%��I���46 �t.Xd�8��؝�6W�()S3��Ğ��P��ݲ�́<m��GƮj:љ+��j�[:�\��*��d�ȼ�ƃA����2K�B�H�B��i�\+P����\6��Qk�H?_	�8�k�����q#�ÃM�ӡ�;T���')����#��F����;uy� ��B�۟`�%i��a��w\��#�����hJ˳̂U�ٛ���Tm��#�B\�%�I�2�Px;GF�;�'%�A�䆆b��C��?yL����99=^CDb�G�kC��wJK4�2T;��q5a��o*t���Ea��́<]og:l-��2�1�P�q��8g�q�="����Cb��|jq�)�V��ӷo�������9��B�:yY4�˨���˅¯�y�Uֈ!}�� eqwp�6n�tp3���� d[��! ��� aƥW���6��g����#�>b�����C�tRuا�G�ɑL�w<~V%�%Qu'֯c_��{z�j�n%������.�6�Y�"���'K�E�a�v-O��N��^�4尕AԂ�y �˿g{E(�z/}����c��:� ���z)kTE�I!�Ƭt�^��9�m��p���}�^�zik��`�R���*-��2N?���jH���6�����ߦ��������3�6_��CGV�s��4�e��?Y�p��1���"u�^'���19�}�Po�	�d@(d��4�{X��2������

q�޿�t��4	Dv���i*:K����y�w%O�N�ίڻ�d��x5��2N�~�
��;����OV�k����c��^������`��v`��R
@.VP���,����m�-E�h��6%�Ru�t��m���9Eo���=E0`3�6-.Ŀ�`���e�C��@�3 ;+>д4n��tu�&�����2J,�v�փ��P��̯���[S:jcJa���Q�эF0I?b�aq|���X�=@�G�#�%giv�B9P������*�y�Ú���G~ц�o���.���3\D�_�vs3Y5������!��x�n-�$hk`���.���w��^�ah�T���b��� F��L5��.��Q�߲ܐ����F�׏�w�{�����4B��R&�Rs6g���.�"}(H�
V���53���ٱ�;%�2o���ʬ��a7�7�KWO*�X�Ԫ߿�
ʏAȺPY!FD���> A-�;�y
c��(�?@̉kY���n��F�*9M&�j6���{~}A#�c9>W�2�H���gjD��b$����P��I�m��ұ �k�-OI�\6He���'�I:�^��9Iw��y��1aG	��hAҨ ��Cr�n�--'g�!�����U�ߋX�޶�9o�����b �S�mt��M_�K ��3��YУ�v�����0 �az�0���%�IG�#"׆b��j{����y���\��@��z��Q ���|ӪMV�N��nC�+ �	��=ٮ���K�}mu@h�̛e�57���� �s��'ɂA�Z۲}KV������/֥��DqqKZ������9�Ƨ��I�= ֏�8M����Ep�+I��0�C�W%kt���d;6�@�:evn��L�O����7���#�ۊ�̬���q�H�1����|M}����ԍ3S�����nI�:�$zH �?�^�ͳ����)�	4 �U�l�Gv�fEǥ�)t��9-)B:�����Jǵ�F�f8��Q�$H9�r�A�%6��띫a�
ہ�i[�~7����P<��{��h�E'�t��E�?�ݑ\K{�"k��T�m�0F0�D����e;kjZ�ʃ��r��5��\��b�_~$:���ʠ0�N|OӲ��SW�ɒ��c@�D�_�K�:�2j|ah���,�!�4 ��Ź����- ����$��jB'���0Z���Dֲ+�$�r��='�%�R��ޠP!ˣ�!)�ס'������"y���\j@U?�[Sk��.������^=�����A��9G���^�b��?��,���_�%���8e6��k�Q)�T�5Z#ވn�:vKI�<u�g��)3|JΠN��2]����O~#����|�֟0�}���p���2A��'��緷��x���F�ê&�`�B���8�>�
�X��-��.B6�.0a�\���=�2o)8K�@�; .��<�s������<B�?�n��2¨=rf���
�tk��2ƌ���v��]շ�uTk%�v�n����O����9���.϶z���&�~m)z�8�㏽�K��4�R+�t���2���iy�I�1W��.�y۝卶��a�D	+������grR���E��u�"6R��0���f�-zI���=>�G�or�
�#t /i!�_�m�R3 �D�e�E���T�w�s��?���J�F	�#9������i?�7x-�ڴN�Vw��{�kh��KRE�~��;�	�X�{���F�ƛ��5\`��n˚	��@�WY�j�BЙ^Y#=[����օO]J.�}���<���a��f�Ĭ�;�k�����e̲���Y�2�]�Sп�Ub�X���w]�lД�6������=�-�i��&���_��{�Q�a[�ܐ�����ok�e?7=\�b�}��,����29:据�^a$��d0
������H�ߝ���צY\ce`^N���Rq�J�.�{��	�)L�_�l��4ȱ��mc,��;z�K��aq�6'-@ؼ�hy�s�%Ű,����(��{�$�[��	���H1�����h�gç��~�C��8��cK�[��	����Z��{�9Y{ϋ�W�l��}܀����r�ċ�7������1Z(&Ŏ|0����5RI���"T�5=��A��x)��o�%\Ma�܆!m��PDz�raZC��@<w�Ho�V�[.7h�x&9ƽ[c�55��e�G\L�{�^�w�Z�t�˓�f/�H@��%C��b�1L���ً��@�殻!V-�Y����!>��Ae:@+��KS��Û�Ϟ���@�ik6��韌oյ�℺��iy��ۣ/͐�!�J����?hI&�ʿ�u����wR�J��V~mFwoe$�g;E�?� ���c�[�v�_��9�^[7��5g�
ROa��ә�V�I��7���J�?~B�����TwCU�<�������8H�J�����J�*LBs�qh�g��0s�ܜ������	T���@���A}P+���+���P�-��a*L�v�^H��VO�md�"_���&�p���k�w��8�H��z�=�6MQٜ#�MAO��_����Z�|[�1�VdZ9~����y�
G�e�Q�7HH�sQ3p~]��,��@���h����2G�T�o9X�4$<�O/��ǜ0 ֵ<;�K2l��"��>jn�g�'����Q	�ҽ�ߨmLkPnu ~���%i���~q��{�"�J�R�R����b?���0���̪�-���$�]f��!=��߲/A�:�MCbo�s��L}��}�A��q�9G9O��&�y<�3���sK.����}#�{�����wǧ=�����@oT����U8v[���f�v���m����W|d���Ys�Ծ�Ye�3�4ļa��]̫���rA�[:�\�@1�j�8���@�V_��{�g�ua�E*������d%%�G�����.s%mv"��"�"�I�U���ƕ%/��e�4#߾��W��X8�j{����Dlo(�K�Y7d�\#L�5����E��!u� [$S�oOl)2ӦE�D�m |]�va�a4(����WZ\���oT�	�H׶Wɻ��vc0M�Jߊ��Mo�2����*����bLI)��s��Yk��� ���	����cr��#!�l��'�Lg�>�g�4%P��%x�Q'��=�N>"clNƪ�)���@L>���-���S�1�<ݪ��(�xc�Fb"�B�Q��L�X]H_צ�˳_ϛ�-ӀQ��&�&k�P�r����f����������� v�!�U���s1��V��\-|U���پ��u��{��q-iz5�N���VB����݉D5����f"�/� ��WT[����L�V��(�W���2��e��K#&9_Zgh9��5�x����8�S"�����O�H���!�Sq:]�ю��6[�e����Z��~R\#��C���/���W H��t"|�
�,����o���6�c:R�Zg�yb��I��=A�2i #�M_��8f��5��3X�߂@Qm�)A����.Ǭ糏'<���r�BQw`uF&��S�\�B{&�}"�]��2���,�����d��ݜ或�<f%���F۫f`�9�,{�H����Y�d��v�ï8!���%��7�����%�㡙�'���@%��yciU�J�'����XGb)�s����B����'s�Gl��	o) ~UJǧ��I>}W�[03��L>6����s���y{15�{2?��\���L�?�Ҳ�>m���r�� �4\����{�@�c	0�=6���:dކN�_���gR��3{��N_Eqqߞ�Vm���v��C8�㖤��hr���������%����W��Σ�듉#�+$�}T�5�s��{xW,kYa�Jg!�ka nc���-ڳ��ލ��X	Z�3E�eCE{��WlF6���L33�ձ"1�"��"��e_�s������#�%����Z�1*n4�]D���I��.��^�Y&�q�OF[㤼�!]_����wX��S�S<l�R�P�!�~�_o2��q���`�)Q�'����%�w�z��|\�'M�{1ڣl��V\
#S]��**��u�D�-O4��B�����{�G��`�Z3�Q���;���R���U�ܿD{�K��z��l�M�UƄ%1Q�bb�9����V�I�qd��X��(��f�l'��}�������7��(�|6�S��]j�qV��T�҇��:�������o�H�4�����)�#�����i��Wm�D���~I蕼��O~��sA?�p���N�,�J��*d���=/;"è���t�}Vkn�\^�3�P-Z�On�u����˄t�g=�G6
�4�ǤPQm��K�[��h��>�kf@��� �᭐b��*�w �>�۶������!���a�O":�S���e�t0y�'�2�Q��}2H{t���)Z��r�q�X3g���6�m�C��"��n�p���MV����i5P���-j�`)���� 9�
tj����DA��>�}f��Ƃ��Kޛ�t[�2��;���A�������@y3�����,�V^��B,�P�Q�9�F�tľ]a#�[��u�	�-ƽh�4�s���_�_�DԒ媻r��I��=�h�i�AN���䍍�����d�n�j�?vx֣���87-n��lG2�R��Q�y�[X ���a�s�=����!pT����E���K�6��Ly�)��#��H}+v���TN%�
�6��;Ĉe�)?(�_�Ɠ��s�\�T��<.�:��r_��u@'���ċ3^�<�{6�`Uk�t���!����O+^Z��HR���X�O�Kng1���ע�+0/=�T�21E�sV�^�~R �L�+<��7RUB�тI#���p�OA��dr O�c��%��n6����8b�Ý����a��7>��Q�s�s�ƿ��r���!7^���l:g�?��[�
��
�i&ϑ��kn\;H*I��\���$�J���%��(L�=���G,��j��O͓C�~T̏����B�۴]�]2���~�ݖ��0�g]C�YLd
^�ͭX�w.1�7~^�S��ꦇl������1`��\��2EѦ�F���EPM�/֧McB�	$�Ah����w��3�|�!���Ij����@�R�j����b߯ǭ3m�ŷ7��{����"V�㉓X~���6��1-�Ȥ�u8,oT�	���a��I��iY��q�̈́&N�� �!�[@H".�����Ԯ"E�0�C�� �6|1�@p֛gD�b�i�=w��1����X��5�&�Gц#a������i�$��^	���<��<\[8a��Ţ�'�6��:~#��I5|�
Ve����Y�ZG�	�Q99���?���fU~��l�K �:�/��3dh�|�ce�=��#��㭲�F �{�K��\��i���d��:tܔR�vI�F�X��>���P�۴�6�8�+�t��C���cƲ��=D�;!���� 5���L�*g��~��L�%$�`��<�" ô�3M0�9_>=��X7�S��������W���LA��&���4_��JV�ش��v����P�G�7�&	���wa7.����v���0@"�A�#lN��ĥ�Z�X����OJrWVr�S����iS���z���f��Oϵ*��sXJ�B�p_��p��ʒ�_�������d6��v��p�UZ���i��K�ٻ�JS�π���Xb�m�c����cc�Bם:�y��8�_�8'Ph��'�c{��7�@�7r��Ir^̝#�J��T���ո�m�J{����U���N��r+�2�#B!�LN`���]zrh������7�MTI�5�6��>�c>�[p�m� �v߇!j��6����� �b���F��[���БC���U�!�M�� .�L��n�q����%q�:J����$�W��;j#4��%��l����▬�3$c��gH�D��U���е�@06��%����	���mj�L�q�`+�Y��q0v|h��{�� ��S�)�W�B8@��2����K;DW�{����@,S����ke���?�$��[����p�h�#Hg���T��Kv �F�RQ�:��Y��)z�t���G��Df�J�I���,D��=�sx��n��DM��6om�r�"rT�jK�1U�����B�	kh�j��ֹF=Ny�[�t�j6̭���WxB���8�VL��zU}�q������!(>��La�K��H���L��+�����Y�~��6%V���P�o>�����Gv���R8L��� ���,�B�x;��!ߦƤ�S��:Y@�Ɉ����545����Tn��nU�3)������C��;R�h��c!	m���y��3�H+;Aŀ��f�1Z*����S	i���vk��}�3x	�jY�ժ^�fZ
ܳR�CpT�҈C�&5�mE�́�B��Ʉ�Lb�.���S�ꃂ�~��/�-,ƀ�%����SM]�Qy�������\�Y���#1(��q�ؕ���P]l�i8c�V�q�^������AZ�I�S�U2?��\ګ�dyw%�rd�L�r�`�#�s���g3lP��\�-X���+�����.c¢`e���C3be�7�M;�	��X	�V>�x��Hz����S!:�Jْ�y�:��uٓY�6
�q\�+P�Pf�7��t��EsLKz�-;��[*̠��kK
���(���X�[ �����)	._�x&M�h�b���+�eb �/y�*q:�c�h+���J�(K��~#�!���j�ʗ5<9��;��y���ws�k�MִsE:w���{�����ń�͞�F,�H�}��A	��x6s�p1|�����2����@���c��7�詡�� ��=�U�-$���~0��k���I�@X���5"yQ�r�n'�D����>{�(~�N�߸����F3q6ܒ��ݞ�˙��s!�ߢ��=���d�D]�[�ܶ#��Kl�O���>׭~�J���+؜���k1Hb�|\�����I�D����g�k�����_F���Z����+q�3�رi�)�OAW�0��Z�H��mwKRX�^���]-%T�~�w��R��u	�m����#BA����ndа��6p�Ur	�,����W&l����(R$A_ #�v�n?�yB��;��Z,m���^AXnb�����0�=��C�S��cZ����]w#���8�A}dP_�����H�!m50�x����t��w���GH���h��4CS�~)�WF�*��]6X�fQ��wv��d�H�i:⩉��]�t�#,ť�M������Τԝ�P%f؍���8	���Q�E��n9��B��nۆ��������q�&�W���]�� Rv�i��k�3 �Թ�˄A�&�������j>ͮ���3z�Ԕ1�'�J��0X:-7������Tg8&�V ���)̇����$-wy��Yra�yb��[��6 Mח\>���w�vB���R8**^Ձ�|)�DXB��IG�>�kV�*��K+=`7���i$���ayq�D��~c0�6�V5��Nu0>XW��a���)�'b�ܦ\(�D�X�T���_�б���LǕ�Ӡ��e[�,��D(nҢ���$I�P��Y!2�,R��E�grl|��߆��Z�Abq\;�����A_�Ί�b���Zb&Q��sO�u/�
V���G����员��@Dj��A-��d!LwԞ&������!f�Z�\����\%T5ǂl�����7|@���(����@�D$=�q��H0�5z��yR�M�r,y�<)>#�\�Fi:j�_�w6����#K]�TTW��ռ�9�~�k����R_F����͌�\<��ݑ�9vpRTL1E�:@�Q�"�Fꬺ|�TŠ�&l�#k^����Dp
�!�
�lq���I�Lb"К]<�2���d��A��+ɖdM�R��=j�{�טUꈐ�9�̽ٹ}ٻ���|3G��@ҿ��-�����G��n
�U?��GRZ
Æ�˪$�\� }k�{�+بΉ�"��ix���Y0��4��S���ջ�dI�B��X�m�ǵ�3��͈��"���t�
�k;KY+T^@�����T�'T~���zF�Rd�o��+餂��c��J�����o��>G}���#K�(�A�sl��z�Į_9�ߥ�<�A6Eh�ߚ���#��w3{�q�
1ޗ��^��Ƣz*�K��z��z��0�(e���y�ŁRl{��[��|i(hW� w�w�FE��3�C�]d�{��Ol�I0~��ZH��檭�-@ã I~�w��z�x-���NM�51��օA�O{�y�`UUx��Nc#M��,J��{��2�P�ש:����d�]�I��o���'�i6���z���e�}[XGsS�
���Ra�*/��u�K��ַ{�o�+�<5��ށ�@���Mv�`c:��s�c��Q�I��]\^R12_K�����lSW��>��{��
Xyj�|�X?��y��o�L�Z��窷G�����v�m���E���;�q��\�����ݨT_��t-��FX�2�LYdUQ�S��H�)1s��{� �/G�	Z��@�j�!�<ւ����w�;&Զ�fa~T��[�c���8�;+��֕xk6�\mcwp����o�E�umڗ�W$���Gb�0�?����cCo�""�y�VTՋ�.�J:���9�]���eA#p��"9L�DoյP�i�g�d}�bo5�Ű���4���(�x��PÔZ��C������B��!��{��[�::nר2р[�v�4#	̂�G��Tǵ}g��l�e�T�������X��%Ú����2J��L]/\�¥��2�O�T��Z{@���Mn����tܞЗ�NŸ-�,��.W��Ѷ�Ȭw&�Zaƺ3��)���,]篂͍U3�x<���{O�񢙉�L�寉�Ŗ��u��:,�De��v�e}'�XyZI&�OZ��Ӝ�e2�Oԁsu�5=�x�B�N�l�ץx��l<�~�b�#*��J/d�nQx�A�c���ZԪ���M�;�UƂl�*
;�s���-��z�D>H��Q����[��n��`Ð��k����+/wm�At�����;4��G�����i��xSG��ZwB�%N|r{;�W��;iW�*�7r�6�=(�\��Oj{���Rj��n���qy�G����g�q�X��Em(1�H4ʹ���׳-ϴ^V�h��� Ptv����)�K�mn��l?x���7ɣ�\	�ؿ�M�J���H�:���1�b�쁦�9�����)/W�[
����<5
�i?d���r����c�hi�a*�c.0���y&{�IP���uToE�מ�b�C"��.I\�ǈ�Yp>=�V�V�ۻ�����a]Ġ�o= dʏMR��f/@#R��{0��W��B��؈�~�eV`���ll�M/@�����[)�gE��y*%��M�֪�q�J�6�֛4S��S�N'p���*'%8�,�����),j���_g@т.��$�e�`x�"����6���%J:��N���1ӌ[�~Зܻ����?c�E29)�ggu?/>����w
�D�S�cG5;�`tU�������ΰ����RK������q��T�Q|.���
�Z���n&���!��)1x�kJfe�1|��$tn�eqM�?�c}�4�6E��Qb(�h��7ψ�[~uj��O$���G�\�:�.�SrǸ@[��, b�����NR�a{�?���CjSk�n���tH�&*+�';�u�Լ�uW~�	!u�]V }(�R���0�s���d|���\.M��xUϗxK���p���oEz0�(���/�<U�'(!`q GP����b���>c�����eq �=^c�MW���������i�ɒ~�pJ�3t/glY������դ�^��S�РDk���A_'y���xO�Ť����)�k7#7�K��'T�N�
s�/��7+���Q�N���-_�W�cb`&n��$�Kɍ1�"�Vc�MP�w6]�q���񭭩2�*"������E��K~���9Ѽ���~���!��燮(h���&��~�Y�Ai�z+}��F���/��'�<�����6��k~k���W]�i!��?sL�jH����.�߆��&O1k�*�J/Q/�:��+�#ޥ(�S��P����̿��]�jp�i���u��k�2}��9�y`�椺%D<���eߚ+8�[�>�x�!��$��Lb�Bq�ml1sڍ���G��$�XW��'��cf�Ub�c�@	�y|�"[�\�V���Jf\����cXI��|������ot%�Y%n��"A�4��!�A����)�et{��Gl�!mw۱sU�W��|lH>������S��Ck�ؒ�>��)2k���a��V��_p@��i��a�EFdC��b;�����jx�Z�D�f�>�,��XDW��
p�ff�6��JƉ��u�1�����F�ز0�a��fܾ� Xz�|w��m��6�)�;�f�j�]�X��X������'���O=B�Ń6ņ;�4ꖰ �����ձ;�w�ƃeo,j�L��AC:,Xd�ˆ�c�Iǥ�O���}�l����L�{�����iD?�IA.��/�zt�kllNBJ�|6�۲��>5v������U6Xs��C� �Mm(��o>J��a��G�0KW�uĝ\h5M"�����2�;�J�=�{|s�㲣�%y�9�$�6;MbAeX/nm�:����o��v�C���砣|�b��~2=�yQ�{p�ޜ|��g
B�ɖ�S2�L*xK�gc��a5����k۰�Q8>��Q�$��5����� ��X0��1�#�����-G�0_�sq�ƃ���;�1�f�ٹ3Ӽ�ڦ�s�r��$�6%�}xt>L]��"�]�Ϥ�;�h*���y9�թ�C�D��;Y96��PZ����<�A��v�����nUQ�2<$�i��.Z{^(��7�+����6P���_O�F�$������ɒ1�&U����&JQtuXЗ23Y��97���0�f���9��L������)�f�.������2�X�^6@A.+jI����!�>�2qs�n�,K���C𷚓/�
�G��[�	�Ź�,�u@r/�'S�V���-t�v���]'A�V{�<\^S�~��*�����8�ӹK��G�K��Fx^a,(��;CM����;��PJ���2���v���.��д�Gܼ��bPe����6MY ���lIF�Q!P�O��B"���x�Č�8r�Z��`�GJ:�W(	�<�3���A�Y�B�K~5�j-98J�����Z�:l�ѢG��\<BbQ5멭N�;�?���$�*�F�$7��e��ϊ�� ǲ���^ 2�u㖢ȃ)�٤�a�ز��������hj����R��8t+�r��!�1Φس�
�7$X�O�2�f,��󗈉���6�mePXXwf��qBY���cl�#u�h-�7 ܪ�V���m%�Թ�����oT����P6��+903�~b�d2�5LA|O�UHH�.����89sMO��N �>�Ӛ�o�KY���1��L#W����~$x�%����Ӌ������\GW� ����ԍ�Ҙ`��p����2��2���n;���2h����h�o�
���jV�uO>�QL.S�B���ђ߾M��>0�����l�����% �� �T���|�߱���n�o_1�����Ymĥ��e����(EK0+�7��\=io������}EI���j���kܦ�����6�	��_�6��R���;�<w<�T���X|B(��@�!=���e��e���_�C�=��>.�H֟T>3$>N\�c'��=��8򣵗T�]�DJ��J�V��iI]�,綐xxթy�G�֤,G�G"Q�[��u���7� ���2���̉#FA���u����I�[Y S�w��z��#�8��1�(���#�H��P�;�!�Y��xvkd���#M�^����p}C�*��g$H?�YE�\��
��4��?'�ė~��0�ǒ$��7�CUp�}Nۋ����W����lbG���i���^��:OE�wϜM�B�p_I媫�9�<�g�7�֥���A�j�%�o %���0Ik�ĿGl��Y�2��9}�����w��`��'��w@L�'�^��f�;���p���Rϓ��h��Ԏ�-��$77���{?`ܭ�/�����@էQ�,�.[K�ԛs�W�n %�ݦ���Es�����z�Z�x-$(&�%ʛ�N��ɠ'.h�a�;Goɣn9�"e��ֹ�}5�rw���]���W��i$�ְbx[������ө^#c�$�%�^}Y�n�w�O�3j�QU)h`��; X����xM~��p��~\�aN��ܲk���>���_Q��|�����`h7� ��{���'���Q�.��\��e���Pn
���oO+��.܉�ezE���[��k;�ߚ2���`�W���x	���W��[r�@�~/��T���q�
RHq+��\��0
@ $1G/5��:���ꁍ8���I=���
�'��iFP&:^ �s�"�b���b�Z_�+�uU&�`~�Z�S���L;�GS��+��e]�+�j�`	����&��lI����%�ց�U��y/��~��p�!f��0z���"
WQ�U?B?0���I�iAML��< �ҡ����At�\�e�>�V���{`Q/�	�c}��)PFTn�I<���� V_���t����g���pZW��,�ݧK~���9(/�2R�dg>���Y	=��H�p�ޛ76��̵9���#ޫ��@Vݘ���1c��/���0E�L�6��v4�K�|-���؇ɧ+����^�>圥��<�0������j�5	�}�X<��4��{4ǃO{y��W�,����g���N�$��������ǖr��u�t�U�J��;��yw-(�=���߽i��n�Wc,�c�w�m�
����ƫS��'Z��(�;}�����_��S�껙�᧐g"1��1?Y,���r<.�O�^d4�D.��ф�"?C,��&u���c��-_�Mx�����Ga��-<�3aT�:��U��:C<2�����*��l��r��tΐ�.J�G��z��TSŭ��Uf�fP�Cx|��]��6�<�|�I��p����8~a���=er�\Ce͓�:N�d�y��V�A������Aj�Cn�
p��Jbe^51�"yP��-���gb�g؝bt���Pm}2$����"$%Oqr(����)@m��[˳s7GQ�z�~��1	�qLDG�r莦����	E�|6��.���,�_�j<Q�0A}ʟDoyjk�l����D�w5]B^>ؾ�;?|ί�Y�09�)w��5lUQ7j��\��1U��C�=�e ��%3�k <����r�SG�no��QbQ^ZPn{���ci���a0�o�,����D���_�dݍ~Z����Y':x���=��؋�<�i���0�g)V���=l���#(��@�:J�RycS:#��Y�1�=�����j�J-#��Zhh�y+�@�@`
���>�f9�GA����M[��]�b�(��	tC5J'l6��@�G������E)d�9V�V������w϶N%"Us�ez�n��5�f�g
��v��7�_`o�:��P��_w�| DhJ)��uUN�OU�	Y���s�����1Fb�����@ �T>�HI(4�K؊L)Ձ�v�����=��y���#��h/jt����.���#﫝qJQ���S|	7�x_r")Rc?iN��0�M��%�l����5��çWz(Yl�\o#�	;�n(�������̔�}U�K!�k$�]��j���5-�QP|��Z>�F�WyJQ�^�����Z0��1.�(_��v���KQ/�Q'��,bg}�a@���!Z�;q�w��G�З\���T��H�����!��҃���nݽ�@�8_�V&=/�G.2�-IX0���ǧ����l��yg��E48�s�������O�xg_�Md�)7�k��2��溊���B������B�B]}�����V��Z��lw���
��_�P��%
�(����4�P/��[��n���Y�)P#����)}����~a����n�IG�W��̕�]�a�u���+��3yӦ���&���k��$�@�z�L����>/�e���3<T⺸w�@�F�+��s$l���yy��峽lj2�\\Χ%��lDo�+�e<��lyћ�ȥӘ� ��p����'Ag����R�����y�A%�� M7Y�T!���:�Q��Ђ�&=���E~������9�v$'E��c�#��@�K_�fO���M���`
{�������L��7{�M���W�7��UV�zΣ�E�7�4�28��[�}�Tq���J�-\ �tc��߷�!{�����6�ɓ��� 칲�d�s 0ar�z�ts^<��eLzݡ���V���6/E��$��7_��Z�2��t��`���v��"Jo/HaQ �ON�\ :�ܨ7]�r�n3� n���8��"h��eC�X*��e�}��bJ{�-c���\{�a�Qh!�%�� �����F�Pg�1�A|�c(��6�T[kV�u��ٟ1�-|ٚ��*�醟�Q��5R4M��$2T,�lȢֈ��
��3I/��ַtE��K�G���M,�d�>0�x�y�i�����R��	�,��7S��3/�B0.(��)�TiC<����[q��I��H����`�#/�t�пA����nlD���Ѩ�E����O��y����5�T�p�vz)����v�Q����N�(������Ŭ�+�Fk�j���e��-��������е�hj���SF�!fd�J}Dׂ�\ެ�w_�ƾqÄ��CU���˫�#0��,��/r#��}V��[6	r�Ӆ%p��g��]Ԩ �n3��ܳ~���ES@.�ê�#�S�i�;:!DK�1zQ`h�Z�_����Q���M��#ͯ�Wɻ����+�Ł�o���8_8�tI��
���X3��k�*^��J(�f_k�o7/�;&��U��%�>5����}B�Q����u_���.p��?!]���q���cS�8�4�K���EoQ�B
1J{mK�"Z��z�.�p��R��{&5q���DZE�h�a���U�g�҆��l�ch�sqz`�1���!n�p�C���m�H�(���0��x�?6U�����5�!{:(���Ӏb�M��9C�^�dp5�(��Øj��G��
��.C��݄c�[ؕ��&�C=�m����Љ��,��NSآd�@Ĝc�����AMK�,�07�އ#�0|�
��\��<��0
�a�@�D�� M��	.�t3Fx.��Q�xλ*��A��/w����hhX\����sg�v����j$�.�,%b���(���p�:�d(^��J�jT�IE��Z�c٭���	-xL�Tg�*ӣ�0�]� $���lD�"MG�_��̮8��0���J���?��0�:j�����h�`�a��8�3���2�5�Xm+ֽW��0���t�hk��k��ŧ�x!����c��Ƿ��i�ו�X�8n�o�-�eZ�v�P��V~zA��k㼤ff�S����_K����O����TPc-<�M[����9t�E�mm�<Y��CV���`\� !��Y��!�R��H(=�Hjdvۻ7�(�+�_Ӎ���y�Xpe}uiӰǋ���U|���m�g��N�c/zv��-W4,�kх�ng���TBt��&��'���DS���2�;t����ŪۅX�UZ�,UÏ��c�p��ޒ�R���h���EB/�n�'�N�l2}2�:g')�:�	�4����1�ֹ�%cɚzv��-��@�X�bQ�j�w�G�-�Ct��cL)��k��p��r���VN��ã\P���&��|��#u�"9������*���f��6�c�U�5z-)��=�W?s93cTo���y�JHx���v���z ��o�	�&����>�Ӧ)w�H���ՎY��:+D��Ʃ��N�;���B�YA��7���}7Zٌy��Ȁ�]�Ι"�&R
����w㷥 ��}x�_�ZE�X��q+)��M�V�'��}�?!*��5�|i�gL�5�Gb+��|'�:V�%���� K��vXM���;����5�������N��Ǿ�&�=V�+/[��H&�@[J*��.�]A��״3�A���nX�&��iy $�\|�����Ԙ���J\�ӂ��-?U��<���b����+ɶn�<|D�إ2uvPxQ��o���zE�FSct��@�z������G7����C�������W��bOF:a.�<p|�r�
D�R���N��GWpM���K�̪�x����h੣�d�Ғ��F֌��n��?�{�r7�Mڊ����·�	Q���`��m����83�^��LZG������Z�D��������0Hʩ��S%j{�s	)�y�)OÎ$�nƂq?��`�7�&�'/�GK�H�wk�H�A�M=��aS�\��ǻƩ�]IZ�l��}Y>r�.�[Ň�M��[��+S8�Y�w����A�4��g�d�ѣ��ߨ�����i��0���L�,VA�Eecj!��v�6��eڀ}��_��ޝ�m])�\p*�,�j����xJ,�lh�� ׄ��ͱ�Ƭ$�z��7��ZJ�=�%�]?�0�5�G� �r��)䛹�?ģ���a������+ul�Y�;�u4?=��.x_��p�s�-�.Ũ" �8�51�F����8V�߷�%w�q��������]� ٰ��Q�c��J�4h1�����X��s٪�4B��\�i�J���6
*�p����;����v�I��[���4�r�Q���Jp��U�Ce��A؁�pQ�x&LI���Ut�
V0+�dG��0�J�!�ZW4���BD�'hDɅD��y��T���J��fS3�pvСBS*^����6D�?׮�\Ge�q�Iµ�嚑���2p@�	��[��[�Q3#���A���az����S��jz�r�+2(f|���0Q����"����R�X�۔��suj
Y��^/�co:��G��B6�O�p�Qlߛ�~@d%�w�>(�~s�J;>��|�x[�/�~�,��v6�tHOQ$R��~���n��g��~��:WCf?�r�m0a+�$�������NN�Pen��Z��vmP�P���k���1{;pwU���(n�_̳I{<��@sE���Ί�*x��-7��I�c��-���>�)�c�id���L�т?سt8��� �l��=��܈����b�d��_<z�b:)��C6���䬰�@X��V��.��Is��%3r˹]R�߮v����)�Nn�F�#���@S�pqVYZ��U(1E�]�CZ��$z����ڜW�t��X�ƕ�M�'��?R!%�����C�w~���a<#�p�r�H;`��ܒ3z�Frl��-y����$��n%��<H�p����f$@sX�(�Np"�la	�#$�z�����*;�4���{�@��,>�&N��jGP^Hh�������\��~KGMMV�2(�:�)f��Ⳡ�[ۛ�Ï�5̴��)OC���C_�w��/N����&�Ϡ"Aq�i.�`q;_�x��]��}�ar���1w����TW��[_�a��,�ɸ8��-�U�f��:��.���J�������9�+5$���Pq�K؆��.��;1���*
��3�Ữ��F�-ޠ�ϊF_8JD�C��������f�6Y���ʭ/��{����5��,LĄgMBO��"����_l���R�I?<{��*������}+S\ \7W������9�� �P�}�B� ��{��#PҾ��Bǔ5��Q�RJ�(6A��Q �b~�
�/3<{?����	�w�ڰ�Ϫ�o5�(X��$�&�KsM�1�Ґ>��`Y����(���UCP�u%��Q�[����@πp�K�c��j���g�.�^���EA0W���C��,Q�zgXf�<<U:'�'�D�O���)���(�T����Ǆ���+�_Oj@�9��W�ܟō���4�����.���)Q�+� ]��*lS5�=�L{��j�"a�搤X7�˲�I���QY��]{����GP ��y����?C�@����/��a@(~C���歇��GA�T"��$g,_;����(�+�%�Ƃ�<���϶���ЏCM�+໋	Z\;?���=»�����j�V�.��@�&kŽ�k���m�-3���M�΃�R(�em�a�Ϥ�U��U����Z�u� �q(������tDσ��,�X�d���'�K�߻*��A~��� �H��1��4Wku�� ���V��U,���U1���ٜ�*ݑ�o�C��.Z�[V�L4�~##����ަ��%��y��ElH6�Z�''88p�GϿA�<7��l;8|�-�nr�~ k_��`p�s��~�Ei�⏱(C�A��>d�{�ID�;`W��y1�^��j9��s�ޤ�E i�T@���u�*3�E/�br�l?�� ���=E>� �/H���URVt�@����DT"���)|�'fY���-�UhJ♻�d/���:C���"��K���?�����F�[��_&���bI/JG׻�RE�0;���Ŋ�!�jYI�����#\`���X����G�m5DR�cD���!�	qE��A+�
d^�|�n��Ϊ�ï+P�>jO�du���gPQv���Y��2&+��c��4u��G��4�PM��f�	���p�o��Ți�i���q��w���Wq��Y[ˀ��7�����+�7�	��ˇ^��!�?~0b��j�m�~]���=���/߲�g��i�:E�W2x>����"��M_��,��PP^��S�g`���C|����]�g-�f�6A��vDv���0��%�X����G9
V�p��$�09IÎ���
~AGEZ��R�u1&8\��l�9493�}|;7!2��h,���p�yz걔�A�tf�}�]scf�5�V|�5s���҆3Z�- �~��� P9x+�U��&�������s��Ε=�����t�$���z�c_cC޺��g�����[�(v+~�����v��������^�P���r~F�?�?�&�m�$3H�2�ꚿɾht`�A��^��P�[i~
���#Y�$������r�Ń��)��;6���|/�ʻ�����:ݳz��I�:�s[QW�^WFu�������x~M`���mRcoH?�F�̩6vxbH/�F��d>I���+��|�'��EX-��x�+�#��]�7�ƪ�\�M�ٳ?�uˮB\C�d��s������2?��L��@^��Ƃx]QF"QK�?m����ɯ�t��w5� ��9�c#��ծ���<h��<�,����uWFk~��HBJbj����z��?�_�4`D轜S&�m�^h�^�I(1��D	6U���f��������g9�C$�|����<И���ٗ�s�-�f�>�5����������i��UKҜ{����p��=���M�t:N��8aM�:B�gM�s���7T0��9�`�f�f�;�҄7������Ϳai��nzt|��&�7�&{P�l��!�5!�˚^q�*��U@r�(Sy�n0��
n@��fT&���c����Sz�c�ߢpOI���puҫ=���fV䦹"4�[уC �F$h��f��ݤ��'��k�k3��iJ|�I�ߋ�����(���w5H�f� }���1�1H�;W��[�?:�<�OĦ#���m�PM]8p��uT`��
�d�}��:f������A)���{��J��iy�ZvK��WN�<Ay�&TE�Y����A�(�݀�XAE�-��F��0����Rsݦ_S�*e��у\&�1��)�u
�[1h,�<HP���&X̗�$ P�E�ZDC��#��}4��`!W����YϷ���Q=Z��[����:G�7�t�9q�3�Dȟ��֙��?T_6�֤	�*�y�kk�����C��A)�4�rs�j~"�W�u� Md�p���b'���zX��������t
އ�� �h�L�u��G[��©}خ2�9�8��mI� ��:G���(������ �ML��1�g6����e��D4Dp<�G}LJf���Y��Y�&P�XV>as�Us���~�'�I�JW����y1��A�%]��ݙ &���vӗ�\萉����S�2���a6oנp��;��<�S����i;���'�{D��T]1򱹥��)#\�Ԡ�4�=V0iDw�L����C�8��x�xU-�?��`&���:q\�N��ǎ�G��t�]�?T���wֿy�v�ݜ(A��%����l$N��w�[�i.�s�0���3�n!T,�,�%XzuÕW{�υ]7n���\ޘٸy�'��<я���Mq���Z{Ѫpi&�Ǆ�d�4;®���3��tZ�>�zǔ�Rګ��3�5�?�9zB�x�G�_Y�E��O�f����;\]�Zv��7���(�	�<�&gۺl�5���mC}Yb����'� ��� ��2L͈#Yoy}�;�%r���0��;�s��Ŷ��}���s!���H��5@�����lE�� ����g���5�*Ўpހ�zZ Y�\�׃X~ 	c��xI�#�(�	2��������	�G��5U )zJ77���Q��?���{����xr�q�W��vo�j�f~�'ըS�#V�\}�o�7>���b�Q�d!��L��A����7�VJ`�.<�x!��ͭd�^�9X��!����Y2Y
SJ�e���X�VD:�I�q�J9�[��[���T�b��U;G�FyK&�W��s�q��Va��F��!8��<ᤐ������&մ�Q��]1�y ��T��R���](�}m	�\����^�-ɚ[h�~ ]u�ex;Z�d�{�]��b�\g �7�%�����_{7W4��
x����+�}$}��e����F�&�d*��]�X��LOk�FvN�QH�_��|���n�i����2"�5�[�����.��<�G(vl�Ag`��j�S�0��f�pl�B2V�_Ӽ��0���y�o��A��̱^�̕6�Ch{a�I�c����w/$ 	+U��cfD�o��q+ET�KT\h��$#V��V�֯W�1�>EN�r����%2�J�#��u���
Řݠ����?wcV��A�/BQ_�qy2�Q��Ƅ������ו����Tfh����3�F/�H�z�B�Sv<U�]�R���6�4�_"IX��b� n���&áP���ȽR�<�V�l��bm}
��0z�`�e
������~��G�.һ!#��V@SZ��;��(r���m��805}v>����/]T���aކd\�7٦}֡:�ր�s�}w�:�_���%�cT�L�_��ug��Z�S����������c��2@�iE_��RO0�cS'3x�bYJ{~��;������Ai��8�3�T��� �c�L�s+�C�~��ɳۉ~ Ӫ4��q��t1��l��9y�-? !�c��^��G~��=A!4ު���[�ʮm]%��G�y�D��	g���*�WY���d�'ɜ�0 ����K�i���W̋DkϮ��o�F��m�d�|y�eS���4���E��3�E�&oS�K��#��PS��^������-pS�u.A�/&������2�7�AE�G]��!�=,:��/���Jx<aL��Ke��L�(A�O?\q��y_��|i��k$���A��ֽ����B4��%���3:ft�Lv�X˧�`�Ůw����gHHb"�4��Xͻ,=��LY��IIŴ0��U��?�J��F�e3Ő�_��P��zf�5W�+��qd�p�7]d��<K�i�Tdj�m=x4{���J��O����i�e�s_R����P��ht�QF��8��xf b2ݴq�s;�&WA�G剪h�fd,����Se�H�&��}�C�M\b6.�iV��BlA�#/Fw�@Qؾ����Ɇ���aU6�.�����.I�1]kI�1nU���-���o�W/�����3�*��J����9H'����߀��0����������Z֊L4�
,x����^�4f8�f���Hms��$�j�P���|���>`�d6�)�h�F�8�`Y�IU��¢�������
�[S��� Kj���K�uGه��?RO�E��J�I�Mt�����v`I��|���~*��N�8��/�/�@"��
�3|.5��.#A��f����`ܚ��	�tQ�C�U�Ygس6kg���`(-bA?�ܟ!���>�Y3U4iX�D��;��b�6sݝC_P�����r�H�[~�0�r�/�
��3��鿡�Q�C��<���Iv��B����:�Vk(O�u��+���ay�����r�l�)Ie�|�*�o��� D�)��ؽ�)Ҳd�yjǅ�h��Qn	(q�
1�U΂�@�2��nnHF;e�S+�?�6�xpj�&�Ѵf���b���>������ā8�:�5�i��5��Q1�9�^����_s}���I�%���M$]:\�Z���DCRit��C����3��伭I5��JvŲ��k�d-e_��}�pN�8/�����4����-��"qp��|�L8�Z��q['� �J)������8\Nd�,��������9��]
�#m�Y�0�v߶��������ႮM�sK�7r*~���H�MБ��%�`	��ؓ�1�֣�+ʄ�a3�[:�'%l[�F��m`��!9���U�����7o
n���Y��Cۍ[y�W6M@{��m_��s:�����*�&V��L�T��Z�������j�aÁ���U�qϟ�DR3�PI��E��KI��泵p��#��ᣦ�\�eA2v�Xxm��a�>���y<���M�<�(�fͽE	59�G&}"�,�:�1k/c7�T<���'`g�S�ęJ�s���W��%(?Z�+c*�ϳ�֥�m7xHFu� �3�[��0��M�ȇ�O��A�=K [��Jt����T����7����ÆY������5΢1�ӹ5*M�j���k�ʅ�E/�)VK�~��j��XY0��խK6k����"-�'@��nJޕ�Jٱq�*^�&~/���(��ӓif�3��^�D^��$`O���Cp `Í�	J�#;tqޚ�ť�^�%)��$��'��Y��]x�5�+���$0�
�5!���_��{��6�i��Q����3���s�E���_�K�-��L;�o$9��1s�3�gv���x���D;�Zj&B�o��ɾ�A��w0��)���>���JƲ7ے�$���l�3��f�c.�J��;��O&C��T�؟>UG�B�ֆoYHZ��%�;��փ�O� �,� �@&��f�z��g:�Vn�yӃ��_��Tn$&3$T{�)%�2�g ncd�x��&p�q麩�-Uj+l��<�b���s�0ml	{�JG�ϰ��;�:�f�@��=�0ӎ$����'ۈ7�_�>������=���$��ç�\� �|L�0'�?��Զ%w�>#P�̝�&h�^��Ҿ-��F�nM)T
�>`~�7M�� 0 O�A�ë�7��c�ڶ�ͨ5+��8'��˿8�=r�����o>�}QX3�����Y��o]��}�`0r�mhRc�wG�:{B�ܺ#�$�� &�T�#�c=�h��Y�])�F<�<WR	��2ttW��o���ڦ��� :�W�3�6�`+��_��~�R�~+SHA���J��x��(����Փ��x�@8��7��w� �M}UXjo�j4��}xQǩRK�����I�;+3���H��o�_s	��hA��/at�՟�vۉ%�#��Q1���BO�!�Iӟ3��՗9�9L�pRv���ћ*�j������E�Rޘ��N��6���踆;0���t�]�J���>JK"���*����[�g����,��D�v�s+uNPJ<�v`q����9g�N����ec��US���o�F��'�b�m˾6�b�Rꭵ)����ˎ��ŗa?#Ӏ�WsMё@#
�B�}��˚E'���z���eC���k��y^/>������	8�l94g����O��Y�O+t��Ž�X��qMt���fXMk�ȑ6]/fsJ�V�Q��)t���E�X7�@E�R �`p>񽖯��Ò���?l���*ޘ\*<�qP��6lXi����G&F���k6���G��T�~S��t�0ۘ��;�!��`�R��#�V ����
%4���Cx��Z�Md�o�@p�K��Y�=�!Vo=�X�ko�;V���>fo��TL�o�j���Јb�b���܃U�MV(Lf �d��L�z���־�w�(R�&o���`�����xֲ��XB9L�e
a�qcٗ�X�8�3��7q��p�o�<+U�V�K�Я�JP'��P�+�3����4e�$j���(]����n��ӏ�و�? ^��8��9��f���k/G�#����Ƌ	nu=ЗB�T��`o_%�c�%�B紂R�+<`�b����dV��$���]V(��J��9���>v�T�ϜQ�:�� �V`��}^>ݲ�ʄ����Ɉ<�ԥ�����DVg���MhZ�VY����O-��
�0[��j�e
{������&OƗn�r� ?�\ReFl`��=�I	�� �b�ap~R:İ	I�d��o��Ѕ���8[��.gT�N|����u<�����~c���^0�+?�)|��{������۲ռ��H�\0�ٳ��7��I�:Q%914��w���]���]�Ӥ�~%�'�Q��N�,�Ӻ��z0s}�r��N5s/��V
�����]8�QaI������M2�I ��	�P�FS�;��������n�������e����h��@;�WT�Ƈku] �����m|rs�/�N�Z~�aT� U�O�zh_z��|1,G*�oVm�A�T�Nd�%S�PXc�8E����T��Y��F�D�ʔZt����$�i��z$"L�7���|�Q�[	UQ�z��B8%�� ���m�9�����X3��t��3\~�8��I���f�ڢe �8���'����#Ʃ0-���jY�Qs]¯��F��C��HX����xH�O��ۋD��Z�U�׆�����~H�l��A,c�I���;7�����f&�T����C�n*�EQ��r���'Y*_/x��J9���
*+���hdTn�"ѫ�kwT�M�q==�
I�|�m�����)�/�O�=o\87bĘ���z�{鄡ʥ���\�����ZWQm��w��ݽ��>�3�rL� ϥ>�@�Ǘ(�Φ�5ѓ㺋����-w��M�>������\[W����@<f���81~���࿕G=��f!��h�7<6h�{sM�'��=c���E�7�U��c6wD��~ZHt%�"o+59yY���]f!�c��D����D�6I{�_�@�yD�w�[/�_$�OK����PP�a����
=b?�U�/���7:i���93L��b3.B)$]tʐ���:�����Y�� �=�}O�k[G��q��.{ļ�U�{l��/�c
�*�ZGI\)$Ǔ��Ay��LQ}����D����1q�ST��ǑB΋�-p���B��E��8J�J��˸M�� �x8�a�����X��ʃ���;V7{�����9�6��ҫ��5��s'"{�2�3�sw��I�Q)4�z�q�aĬU=����"bη��V��Fi��K�C������G�B����8P���#n觬�$�q���2��}%��4��R�G�)�_�7'�;{�pg	�X)�N�������M�׸���ߤ.H����Ӷ]㮒�	�]*31������4ߛ<�d�e$cn߆v�#z6�����+�&>�p�QG-R�wiJ��6�8`�3١KE�:�J��T��9�~w
X�2�O�\3��o��D��"i�[�lq�'p�iSr����9����9�_㋪�z�i�����L��]E�~7�ˤϐ<�6x%�������vܧ�'I9�u�����
][��Z�P��0�����x�(�����풌 ���ޱ��L�9�ߏ��>hld�ė�=n�a.���b�yBp���W�ӈ�k���9�6~�b)L$���zgD�mG.��y��%	Ջǆx1HG�A5�����j�����#�f�&q��1����w�2�_�`���^�M��W:��.�/�మhd0eR���?S����.<�`���nm���6� X�"=��3/}��2���Ƭ�V8G��"�9�hN�U짴G�/ݞ��C��]��NqN���U�w?\�i$�#B3�l��[W�9F�ˠSl*�Jг�^!��C�Jz��bx^��2�	:m(=�{v?7����qU#�HF��N
w?��%��ҞGV��	u'
]-�S�p'�OF�þ�����ổ���ɥ����b�[��,�쮽��5g�G� ���%.�嫀����W����n��I�o����ӦuL�R��_(��]�Bi��{2%H2b��f�l�.�ֶ=v��ٓZB6I��z�1��t;U^��b������OB>�r����X.�:��Q����ۉ�?9����mSY��Q��56�O�>jIB_ę% ���%�l���&($� �����U��c�JY�p7Y�D"�BAu�8��yy�B�Ж��	�9�"ٌ��U|X��Cj���;�p@����8?��ϽI��yu�<T��m��a��w��{6��<���6�Q��t�|�U}�=��X���G�'���gQ���d#40>��}nQ�c;5*����&�PoZ�-3�Ϲ�:u��@�"T�\d�O�&��xKz��4>�Vg�3�>S��Y:Ý�� �1b?,	����O��Ǜ��}���MC�k�<�bt� ��_<���5�B�7�P�|�P�G�7g4���fR��TT� ڰ�!��'�F	Rݠ���/N���2j�n~�h�6)�]��,}�A� �0���8ß�Y�T���	,>e�c�,&�m��5�q��> ���r�5:C���m�
+��5�"n��Ӵ��;>՟琔���1�������t�D[�؜pO��=����=���zf�R�֛��:�/��l��� ���<��C�:MHro�G���ir�^�̡B����'��ebX�~��4#�Yqe���ahM1A�YsL@0�u�̭���X��F�g�Х�$r�r��)c�o�'j��X4f�W��V"�����+�A؇���;)N��KwJ�ѪbI�Z�(��m}�K�U�N��q$��<{EI��1\�<��%��UOۍ#vz��P���Qi�ph�:'��X|��A�~��*.�����M�r��%7�C.����f̆�S�Iac�xB����@�P&�	G�ю��4v�,��V����|v�࠻ X������F)U��Hsò|Qf�N�j��!�J�ǅܓ�3p�hI/aW?��c�$����iV���Ysi2��˃x�ٺg\�i�*"��
rۿ$��b�Ը���yE�h�pD�_�@Z���b {U�1�Å�����ן�e�KZō����C��5P��8R�̰�	u᭰��$�Ƅ�^�H�����!n�:3R�V�]\p�lx��>�_��	�:��[%�j���P����4����yk
��aS�Q�UY{\(�`�h�_q��+4��8rv]�V�r�mC�$�?�S�i�}芰̯�W�O�����qR�^�L�$��~n�g���S5y��-D&���&��@�/ ���֡��Y�2F�>o�T���}��jla*��1ɪʉa�Z�������+�=��|���g*"/pX�af�&H�Lw����?D��/mR�\���n.a�r�b��j�!��>Q�n0�k^��̨�=Z��^V�!�am#�э�;Cep	�_�|D��p��jb>��<eš(@���WxE���I�2*,�_�J���AH���F�W&!;Ze�[�ÖW5�BD/Й���=����~�[o�Az3m�6hH����e���#'�x꣼6�JQ�’1*��Q� t�~@F�1Tm��ji�h�kL4�#}RL�+l�1!�[��H9>�ȹr�f���r���k>�|;J�2�/m�3��[wԫ��n����N��ʹ�#6�D�K�HKuT�8�t߹�/�DawY(�:��`��溰�[��٧���#iA�r�/�_��i�ro��h�!�œm@
G�O�,׻]���u9G'��V�)wT��g�����ɩ������o[���?��jb�i�(�k�7����&q��^�Z{q<L�ԣq���u��H�n� G��tΙkٶX<͢�1y`�ʕ�^�H0�}J��ﯸc5���e���w�a����s7�33R�c�5/���9R�ʼ%uk����4r* �I]xA���2M��(�#Y网��P��2t�˖�O�0ȕ;N���L$"�H��6v�YߧDT����S�щgk1k�ˇ����FĽ��.�@6&���m�N_�rE�\���=\b���=@@��,�@)a�S�[�Z�ω/e�A��� ����;Uލ4�C��C��Z�{����X����d���c�_O�PA���E/�=�,����f,����н&0 c�p
��מ�>FP��H��UE��c�gO9GP�4B*eE�ez�R���-z�f�	M��)+���
����_�b��C�g9%+�Ktc��P��k�y<�Be�&�8o'�"CLؙΰD�u�����Qf�}�R'��O���
�|���	N�n�;�.ǡ�����C�s���i��P��gPo�,�Īm����a! ���"��=�Z�(<����D3�`�Ű��D�)=�9&C�����ݾǬ?���jߐ��}�SX�?�J��V���/�0\A��BAEL�[�y��'�*�A����e�C���imX�^��ur|��9"�_^5 ~��8���WN�xB,
�h�ӏ�P�q�J���Qi,#�[0�l���"zaJ�>�H��W9��IY�&o�(�W,���m{ƃ*�H�2g�	���%���6�^���rM.�}#�3�R���\1N���*4�Z_qW����g;��e�Nnw��E9��>G���;���O��D���D����ۋ!�+���fZ	q5đ���@� �6��k#8�����VE�%A�{�7��W�Q��g�	�˶�C��,*��mK��Φdn1c^-���ܒ�\�g{�.��89%Uuח��O������fs���K�ݐ�Ғ"wm�j�Uq&���wĘ8������AG��ĎSmgE'�7��\)6d�(ՙs��cg�L�ث4�����~�h�l��3���pO�-y��(����#s��3}z �����v��%�U��]pF"0J�Bm\v�^��ݔ�c�.��%��0n(����}	>�"D��ćvl�R���a�Ao�����yi�*H�;9���L�Mh�R��f�=i�k��A,uQ1��
+.����iFH�`��ѣ���1ת;�Y�6ঃ��Fz��ߜ~�0�������յ�WQ�(�d�hf�!
Ⱥ���M��k���)�d������_4z`̍�	��sUMc>�IeחR��W�5,	@�$�d?�=F���l���I�dk�;t�dl�-��P��S��I�b$�j2�P��{���i��iQ�z��)�A�Iox�a�yFA7�$�V�O_�"�)�ޒ5��J��9��X�&k���86"�ψ�[2a�_�ϗ0Dv�MfY�KB�0��u�+PU(�sl����YY���w��������1iD]�T���ƒEF��<�_��e�c2L�>o}������;���:�d	�N/�� a�
��	�����<�;�r�e�w�ٸa�I��ǭ-#`��pl�����r̀��Bv��@mA���M����������"�F2C�� �li$�pc$J���[��
�	�����%���}�2�\��ο؆��ʁ��
 ª�_�1������vW{���/i����	H�u犀�C����~\.�bV$�#�!���Z$�Ȃ��d�2���.������V��AYp[ɣ���;��@h�Dܺ���,�)�|Y�!4�@����+���E&���=x4��I����A~��iN�����A�J6��+je�"�94��#\��$Xxb �6ų]},ȧL���o������2��GF�1x�م�pŨ��N�q�
����s�p���[o�L/��V����~�ea����nd[���"ij�.�T�=z�y�>B]B_B�u�	5����Em�b��RX�_#yi���� Y)�rO�����d�u���x�e��u�L#�r_o_�d[u>ZJ.�pbWjy���B�Pմ,����X���p�D��F���I��ӭo����p��+ ��@8�sC]��ꟄQzWr*�ְ�����f"%��@?�J��/��-v1nM�n�F��Y�Jbco�D"�^�g���K�E��&C�.VZ75��6k���7���#���7�S��RӂF����Ʌp���b�����J��4ő����1p���h.mj�lټO����5���@�W���
�v�Ҳ��ƀ��ߪ{y���%SwG���6(�H��+Եm��y,Gx�?N@5Q ��+��|17��� ��3y�re2��7��{?��Ax�Y�{��i��+KpƋ�B{H��%�)ޭ�U^�� �Kӳ)(�
�:]��)AU?��V1�xr���M����n�t}, w��X8�;�ӱ��ï��)��G|�3�Y�f�$?��i���8�����z���NZ��R؂J�6t�]�L�F.��!e;�s�֘����f2��y�R�@������y�".?/��r�B�QK_�a=���n��eR澫�;ͬ���U��y�sM����:��?�$�Ʌ���ĕ5��#�`��+k��s��_���G�㘊2�6�ֶ� �(N��`���7̫�1����k΃1� QH����z���G����__�=U��}�҆ZŞ�
B)�"A5e��-�!%_VYM�j_("A��ԥ矓�̗&��V����~R\��z귑i��h����P�7�a�b�=�;=�E	ȇ�X�`uN�B�(�J:o�(�H��ү���|E] f��rٞQ=0��?Ax�*J�?3�\��ci�Y��B3��g�?1�=��hϠ���q�=������TUi�(�?Q*YH(�ZX��!-U�͙(ǭ-�`;jy+�2���F%�S̷X$�9�5c��M>S�B��}�ݻ�b��|\��!*�7^��� .m�L�����TN7��� ��D��P�l�����w,ET�˰��;N�1��{�Zct�Ѩ$�ŕ%)�>ׯ��7�8Q��P����b_f�<����HCu�<˔,���~󒪱P�J�lw}�t'��w!%k����$�?2��a�ؕ�ɢ�-`s%iP۳,��q:o�!�F���j��Ï�SA��]��Oi�W0{������y��W�S^�,��^��J^�ޝ��y��I� ���C'��Qt����nˇ�\��}�l�C�a��Br�>�x�zO,0���jUa���fN��i�5�bzS��& V��֋�u2eƾ�o�&���ښo_�y���B���4
��Nhm&{\5�[�q�Tֆ<mu�W��d�YVm��]vnN�
�q�H\�Sc:��)� ���HS�@� �A77�=AǏ_
F�R�3��(䷶9[����p���/��(�cƼQ�ŕ�S�X�V���o�������dB��4kd�t��ǐ|�߫�E�6��TE@j�h�n�1L���M�m�g�j��L��1�|�c����fvH��� ��{sl��2L,��X=��h8��� ��ʓ�B쪖PH�M�&�dB�8fxB2�"۬iʵ�����!b���S��.���4HT{��g���Q�lH��y�z�vu����o�8c��D�E��=�(�o�*��NG:x~��E3?ti`g����9�I�,@�:�Lť�H2d$���m�F'?����IШ���}�xA\�+n�m'|e���r=�{Zc۟�o���!������7��݌0������4n0g�o��=�@3\94"���{E���v>�o�q
�τ~�ZSnG��p�����G]����� ��,&�İ��7gOxFf�L�r�z�,2f�K��JKa��6��D�?۴��@3��#�e�p�"���C�BZ��~	�e���o���N�	�~��[��ww<x��Kg�	]m�ϋʸ.I\>����"u�I����	$�T�x��t��6���]�������h�bj�$+l0*���aD$3�'���+B�����{?�W��v��AQ��h�o7� M�G��3����(��
�p�b���s�B��c߯�-�{��R�O��#A�2�D)��fW-��c#��^�\y���om٠yݟ�.А�-h�%��_>�B}MW.~#P�Z�$�jaW�>x�)�n��Q��Mw�|1�@�L.���vo�P����-ƶ�^�)�y�Ggy"�,�irN��9^�V��e�N����s�8``�� �d���l�D���w)�3O��;ZeFH�_����b�H�m�V{�!��)v+�,�8��ඪ^,E/�e�^fP��2ͮ�}��h����q��DU����~�=��c:��Gz����5Z�Vt�to�����_J���RH��cU=�:����f�/�-�v���+�YP����p������܉��[�x?�Ν���3�>j�)�|�k��X��ĕeSG�T.����Cq�Zku>i��!q;v�w�=C����7�_��c毃 ?;C��^(���/�{[��X���q����ܞ*֊���we�g$`��@�{W� �kh���١�%�e��?i�B�i2a}ʢ�j���A�͈ ݲ�0�J�98�����q��pٟqg����c� �FK�r�5���LL��}Z'��S���;�o¼"����`O���c�df܎��;Y�o���?�&�z�R�9���,��p��kN,܃��&����)���(��:�P^?ßg}�q3���9C�vȑ�O��+!���e��	���c�k���+R��`�}CX;�V��ШD�c(��,|�;���t�R�X.�9I��`ɐ��<�0���b�*��;��1-KG0Ya'�,>l8��Q�2����� R8�S�O<�W}��#�+Z���N�y�v4}��0X�����|�l/�L@�JSг��GpĀ(]����|ut��|m�O�}0��E��x�!B���p��׬�B(ޡ
RM�4� �N��/jYݫ�a0�)F C������"}�P*PT7߷�1�^G�O~~��IJl@��@(bݛ�
,��oT�=.Ͼ� bc���Z�Ǉ(�	����m���\z�NE=G0?k��W�h�S�r�	ߑ8��W�YUK��c��9�������&$�{�o?O���P�q��آ�`\~�m:hE]*����D��L'9T�Z�q���B{��O%N>����|��;h�i�;0C��V>t����W��rN�������n'��,Z}�f>皹�t�Bmg��rw�e���^�^��#�}�����p9��:�TJ�{&�!�/�%$�Κ�Ca�۱:5I���nw�&��̘�s�,m�Lo+%��v�&�tߦ�S�놢�~�W�T�ov�=��װ�6]]�Ә_� �=H���Z��q=�{>�ƩWp�
�� V��{�}�g��#��#lNLT�t��D��.X��9�D�G�y�H!��'�>)�H�#�Ã�b����j1n~���D��+�a��VaW`��i˘��4J�k��[Wy�d���O�;f2vo��@ם�j��ЖN��n��8�$+(�O|��/�:wxD�OT�7�����h�T ��.P��䒑)>�������S(��(����|����Y>޵�4��d-�'�q~đgɇ1hf�j$�]-�Aڷ�im�t'��L���Wb󧀱�R�A�*�k�hۇT~N�BkB�HL���Z��wh��J���8�L��m��ք����nV�8L
�/��4��+��FEӯ����F2��@)X����M��L�W֧�3e�-f�C-2�Ԣ��׫B��K�-��N)�q��S��'GT��X�ʫ(��	^j�3�ÎDDT�e_��൭x�9^S�4=��ߋ��C��v�ᯨ����ٙ���>���%�@Q�kP�j�����h�:��%�{�h�v|z.�Z�.�&_�e�3 �v]�m���'�y��	h��Y��2)֋Q^ţ���ңg���R\���&�zA�:M"J�:eG�%{��e�3�eϪ^"�� ���޵����6ݘ�rO.K
�����ᬖ}��n�r���r�o�0	�*xO�FSqxhm|G��&�*��&�����f_7��l����B�� ���/xE�XP���[���=�l��DZ�␉>�
I�+JX+_|����/湨�k��?܏� Xw�6�WN�ٔW�+:׿-c�Ђ�(���!�F�I����yК/�c�h
��$���3{̾���@eO����~�!���'��į9��� ����/�W�u�'h=��(� �O�-���.hkZ��G��X0��9)f�r��>Ӱ��ܼ�]�����E�)�"�-|ar?l������ ��M9d�tB�an�t~����y��-��P�܅w7F���UB.��'W�/J�->�)J���;�xR�����	E���p�4�z��1��̫	���i�&yMUx�"���A�ګu����7
�0�&d1�'���p}�����*��v3+t�G�����6����>p��._��e(�2�rZ�|9H�ql���0H����,��t���E�.v� d��`�H�� f�,�&�vV�+����~��^̕1��$+�5ՆX�%��]@Y� �}�㕫�H��R����c$����2EC
������ג��Rا)Q�|V`�k)�E�'F�� Ȅ;(4ъ)]��3j�<A�����,*"L��H�GB��K��Ԅ+���I|��4������'�	8y|�U�;F0�0��X��P������t�Cu!����]��A�
|�1U�	���>���O[0)�_L�w��f�y2�c�B2M����<�攸 ��p��8ä4��߶��p�'��
�^����j9���c0]����%�)��W��
%��ʤ
Z��������)�����LΗ��l���w_1��p��W+��ٕ:�ݪ�	��I�x�*R����������PJ��78�p���?�����������	f���4���o3���� rnOE��lQ�mT�"<Qc!^׸iΙs�f_"�ػ �g�)�ʽ����Q���_M�*1�Zl|���3�c���D�Ք���3'A��y^��']��gr��[T����~���G��Z-Y=�heS���x,�#�������������!�;7e��LbY�A:v��f����GH�&0���+�q
V���c�o?^�b����/�ĸ0H�6�-�AE�'�"�h9��z߄������O$w'�7ylA"���4HK�;cVt
�Q�!U)�i�$\�7f�A�����]��w���2:8^0L�썬����~pd��_�3K�MF5h��E������B��"VhG�?�&��o^LV��
[����W N��6���-���g���_�x���2Y�,p�0��x��}؈�"!ZUS�)�;$�g�w�$9a�P/��;�0��I�;Y�j�z 'B��$��m3�ET��� X���R�6��|�+� >�H	�
X��4\}ϭ�.k�8��ѥ���\�H�6�O	���|嚩Z%��`�&j����IG��-�ƴ��z��B�
2T-�0<�9jߣ&�����E�P�-"a���Ɲ�Z���1��|{%��_��ʺ���$Xn���Z�C]}���� ��}�T��O�]J4��^���X'@΃��p>ǟ�4��]6-hQ,7����HzƘ&5�lf%N��ǸL^?�o�.���v�-������OH�f^���}��3��H&z@�\��c7�{[���8���+�~O7��Y3�%j�L?����d��N��L�j���D�Ǒ8��� |���-�Τ`ӌ��;�BY��b�)Q:��cDAn�JjUR5���&WD��:]�xf 24�c���oM"#V��o��k�9=	�ܽV�&E̿���Z<�N0*�l{����wB_p[�J���Fʭp{gtK1�F�13Nf�f��+��ƹ"��[ܽ�Ԩ�����!V_�S�K��z����19��y�vs/8զ�p)d���\gpq��wY��T���I�r�����TP0��2�u�7����{mLn�5���B �Tw����{/���&!�71�:�ࠊfR�6��+�w�����̴.�?�n��;��P�ɈE!�^{w�D5�X���\������,J���H��wvП����x1�$�Z�Э��x�� h���6�=N�=��P���Rɺ���;,y�bk�no'��:+J�s�?+R>���I�6�kA3���/��L!i����5^�Ǐ9��J0;@E����~�z,�ꔽ�N��d@mb�#oe��8a_�YHQQI\����H�:�Z�|�tr���:"+�+Z_�1�X�I0��S��1;�92A��Z�>�ƶ��l.(��N�~O�n	�l�*7����r�2�Á:5��u�d��d�FH�OMQ�J/3}������лΞ�	;+"�I�S}��z���2ަ�u(c8ZRO3�b�,�ܜ��F�դ_=�2]�.�h�/
f�����X����������<l
e�c	H�����{�xj�2��D[������ի�ս�T]����Hc��y��Dc3>��%����j%��d���Q�X#<͑.����x�9�'�{^ O�wT�/l�Ǘ�or����t�5��]�w�����Ҟw��W��<���5�?CYe���S4��n%�g�J���Ke^P�H�[;n��ʹ�QR7�4ۂ ��R����
��_�d�~UP,��G�F��:������_l^�=���)��N.�k-ۀ�қK���Ǭ�n����~2���
dn��Q�W�ƃ�a>!Zm~�u���#��g�։L��?�m�	��p�o����f6����:H;�L��x	2���H:d��ZR7�3me��Y�Sko"%��M�5�{��B].Y�!t����	99m�ds5���^EVnq�Z#u�X�c���cj"ǭ�\�?��	�G^�;'��kF��t��,.݋��l@�]T���f��+C=��n�WGCh�� g�T"��-;��T]��`�RAVg��zgS��+���������r��.r�Ƽ��H�#��(��t��E����)�,:��� �Q�yB����H������hF]��2���S��`�#��H�s�h�<sL]�����_\�%]%����$�j�4�i0u\f�X/s��҈EfEF���j��c�h7�=���6	1!��4�ˌ�X/$3G��5��%K��/۷MȄ�9%��õ|$�G\�z9��iXBq��<ԣH �%cu|H?�zt\V���ӿ/�0�W0Ό-
#���Tˢ�^@��Y�W�b�����B�3u������b��|���>!Ļ�x预jO-�
��~e@I}��t�J�#�)�&@1\l�����%8��oI��v�� 0~2���8R�@1+���-"�=2�_��4z)���J��Y����a��]���@�[iC�k�HF�/�ؼo`�M��ċ�[���u�*��&L��i�Ɔ�8M
���'xyCw4F�sElm�?������d�h�8c
(�Y�Rg"��2���͍ ?������X+�����#��S]ky�bb�Y!��t�NeC�����B��.I��U|��	̠ �qD��"��&�������M�Z
'R7�����P\H��R:�A�;˲�Q��O�<�ͱ�+�?��~�*@4�q��q_:fe�_!�w"�1<V���C�m�`~2�4�laB<MFeI��B9���H;V����D�o��~S�U;�v<$��[~�d4F}���Q,��Kr{������jrV���p2-g5oLf@c��[�-U�YLJ
'[+`���!�j���Ef;%��P�!6|ᒹ3���>v�@�"3�>��_�,z��ᇯ��ݘ4RM�oD_��-�)��	���l.>}
iE�GSi������m1a߳!���� ��#_�K�J�$m��6��sќֶE*78��S.S_C���0�B�g�*=F�[m�v���7/Ov��j�rpi�yy�J��������Z� N���zuW��.:��>ӦjO�F���h�
�T&�TV;��rL�ݫ���pj���8��j�{��Ta@gab������R���r��,װi��K�V�m������)�bR�C8�Y]�B��^YJ2�=3���J�@jkQ3�0���{y#�����QjC��.,m �%\F��PZb�o�����N%T8���"��3g!5H�hQ�R�n8`1��j�p�3v�6�3	b�� ���C�D!���+�zN���	R�pJ6A�N�K>�5��e�#����UL��&`�p���ȹ`��V�W|0�-p����ڐ@~W�w�I�5��O��BA���/���n,�s�����X4��� p}�?X �? p�! ��ڟoi�R���<�S�/��3>]?�)�o�M(�q�0V���t�?��a5�{z��������%�67͔�_	b-��4Ez�l�1���gʊ�G�8.�<��2 ��EK��ԃ�1VU��_�����~�n �Z�(	8��������};A��x��=�.:��4���&M�	�n��a��O1�亩�wc��U�Q��e;����-�0B��t�����>��Z�]Qڰ���7�Cv��ƁJha�ƌ��V"�)��r؇��K�\޻��ޅ	���98���&ǽM\�
}�=��/з��F��x׷å���!��@�C�%]1���9�F���)��)K��^�ւ������Ŕ!��5Ҥ~� ��N�LmA0�5�kgst�X@���0���?�M
o$$n���T3)\�,	� c���
MҒ�� cdf`���-�$�O���ו`�G��>�K&z�:��S���k�P��fQ�c��'��4�fO"X�_�2Ă� �N*&�B�s���ό�9"EY?4�0�F��O�hy��$Ⱦ����n��i�n� rĤ���HQ����ż�A�C�A,�)H��Ǻۯ��=�!5����y�U��;���냁�
�m�t��t$f�������z�D�eF�Ԇ-�Lߏd�k�1��z�t�&�oO�˗���ɞ�� ��}���mX7� ����8g,#���k��2=�8�s�˺��.l��^��=!����;���X֠*dN�wY�Ǒ�|����D�ݻ=m1pYM��/- sc(:����3,ޱ��_ϵ�ܨ�$��R"���a�n5sG*bZ��(W�����!=��O�bVV�v�-�V� Vu��(
��M�v�g@�-��<��P]���l�	�aX�u��.qz��86�ƕ������t��؃w��r�Ÿ��t��^����Ja|~��x7L�we/�����ob�ic�R:��k7���{R�;��-���
Y�����MQ�cB��#�Ϡl<�)���f��h"��sĻH���:��_u�	�yPT����IO���;�2f[�iu�������^�kU;}���Z��fʱ�i>��[0��^������V��Y{s����H��z��&�JT�R�d	3I̮fS�fe��-���3���KYȶ7�'/r��u�kn�P��#����#,�Z*�X�t���♓�]O�z��QM�Fp�{u��� ��' !����s���4�����:���=�`� �B*n�{M?�L�Ŵ�A�z���e��_��ƈ�=�f֞�_J�mt��q��k��ʙ'�?5*��ͳ-X�cqFf�7n����j�3=V��0��o���-~�kpA>H-n�����,uP_�0�0��L������p%UK�6{��h��uҙ���Ĵ|!*+�Z�?�8�PM����ڈǬa��Ǫ3��(WDX���p�p�ƶ��3�L�A=�����z��t�Oh����L =&����+
�u�ZP-��0�����+	��}���3#\Y�T9���	���+�b)�	��k��3�M��#�<�`��� CA�J�@F��!@��p��s?���'�w��n
N�`0��>��s�(���;���(�%FƏ�s�<Ffux
������L�{uޔ*cޱ$����d�:�wCdN�t���7�{��V��aI�:��O�ؒ����js�N�)��c�5�a��RlM��-�)	�DN[2�H�ZJf���߇�3��:��3���*|.��[���yesY맖���\M1�Z��z�3�j�p�_�Nȁ��S����~Ʀ��Gm�
��h����dl�@�'�`�7��������HaSs\t[�hN8˦�ڥjx;"�7[�<L�㧐�7!�k�\�ȯw�:���s����m��+�Sp! +$�����΍9M�4���w �.[���@��)��	o�h�eLe+<ySW9�9R��Up��u5�.�U|kb'1���c2udx3�<}"�����6�˓�V��b�f����s�uw��;mC��$	��C+*�m7�*��G.�U^�@ւ�]K�T�9o�O�~�O�IM����y��u�����sZ�A6����&zP-�ynz��y!�C�@��1 G\��_V:���ZCz�ٵ�+���?�T\d��'��4闵hzM?#ת��Y�Y�B{Tm�Ǎ�D"oM���f��Y�RFzw�^�������~Ȼ�r�TI�5�Y.��F��e.��\&zֻ� _�r���mI��>�W� �$0`�W��1�#�`������U�!���S����8�'�e1�d��PH&�f_���GM���h'/G(�Ƕ����^$���QO��aY��`F�z�a/@."�gL��"��-��E]Z���=q�
�g*�a1���E{G���~����ۤ(��t�zT����z�3쀶+4IPQO�xs>юlTqq�lF$M�:�ğ)aZ*�U���R�*�}X�j��������+{����$ 
��K8�=*��^3a�~!_JpmH#�ӄ+�f���鱿A'~9tZ�st�z1�n�h��U�۽,�6S�#8:{��Im/����[>�O}N#(�KC���/��0���6����B�O�j��rʜY�{�T��d{�7�s1[|k`�Kj얝j�pLC�����T��G��g�ӷ�ԗ�A����7���b�2toľ@[�]��������KO`�.=�m�^]�h;%Pn������(Ӻ(5����K�|(�+*F.�#���4 ϸ�����;����P<)��G}�`O�2���'f[J<J`�Ι���<����A�s��F�{� �+��-e<{tlS7��f�\<���(���PnV� ��F�J�T�����D#��2��@s�nC��F�5^PQmaܱû
a��?�5�{Cp��Q,���ٷf/���q���
�Nث]MB��;l���BY�S�6R�9��	S�3&Q�q>�RBί9��(��O��FeA�+KQMq3P��0[�#G�)	���O�.��A`=C�/p�7���!/�q�
sPI����l���iP��0�b�:����R��%r/J{b��xRg:<iK؈[�	�`s{7:$^�)��G��S�b�Krg���|��,i���Z�����m�#i��� ��Tٴr�b<��:KP���[ŋ�
��lZɩZ���J� Q��&P�ǥ��+ط�������3
�.n��8`�]D8#}��=Ff^�:*ȤH>"�M�Z���kNW�|��;+I%����Պ�v	-����eT�"��'#8�Ǖk��i�ǹ��|�p����5�S:��v-����%���;���sHGkB�;��X�*���Tk�[o�y��Y�|3��k�VM.ȟ��﮲����rw�KK�=��,_ �	X@)�E%R�ٻi+Z�����5	���dV:rP����
�X�*n��.X�oaU�,1V����.�o�T~WrV#h�f����_ �_KYl:.��P�����<X-	�#F���CqR��Ѳ:��a�4�ց`��ʁ��[X�]o�(o�C��75X�m6��
!�ǳ��:v�´��]��|d�TP��y�A4��;f+o�HZ�L#EIs�Y�^�f2����E\=0˕P���}+)��(�e��;�} �e@�!~�.��^4j�����YK� f��)�$���Yc�l����	�������G"�y��qʮ�N-��y���'\���E��j��t�8Y�&>fΈ�NK�--�8<e���� ��	G���ms�m���n����=P^�YJ�pY�L�H�o�^RK����>:U�  �(v֊l��&��V=�f]O�_�/
�L4�Z�^[A�*���1=R��A��F�\��g�yҍ��G�R�wM���^V�R�\,���z�.Q�W4A�`�����1"���ϤN�h����Y)� H� ; Z�&L�%�����=�� *9�t�j	��	��{�~�kFh3ҽ�yeLZP����Va�+5|6	JFT�sK�5��ت�}�xW��{8鶅���0�9��=�NБq�L!pu��l���ѽ��R�&�DԤ�-�5���řSa��'�
v<�aj�8�4u��G�'=f�BuԃѕH6�Xc�F#B,'~��~�:��ڈ���� NU��!�u�+3��.�AH3e�ĉ5����['�`��v�� ['P��J|�R$Ѭz@�<�C9���'e:&g�^/��b]���A�*��eL�,틢H�ǆJ�,�|�Z�]#�#*7Kf�Y�n�0i,��d�t���_\��*N3o@?4��㶾�иٍm�r��!�����*�=
��P�x��0��ǒ�L�������b4�z�.w�hp��LlU_�`!U�Z�vx]�W_���F�x��t!xs����r�~���?f�I�����(</ �|�`˒�65�K�0Ȓj����{��H��j���'/��B ��7�_:�����S9gM��	²����y9ܣG�ʐe��!��I/I�
�4�9�F&�w�Y6�A�pJ�ܙ���`F/�c�&KB�����#��Ӂsʽ��PhGg��	?o
�k�)�ڂ��X�|��
���m��I�l�9C������i& ��$U��X2զ��K�^� �!�J��8�2P�M{j2�5�Q�eA��3�
]�B<n����&�׻&waFq��{6��tQ����pi#��'�L����{O������H����oX�L�Gl4g���LV{�vW��.�Ϸ�?}�]���7y�
��� �-����N$�O�0̜�]9�����z.���"U%�l�?щ�]!4�N/�ǩHm��\ż@�;�Q�*����'9�$�S|�e�ޡa!ǤƮ���аa��6�.@˃#�|^q��0��f���T:񗷈� �({Q4�a����}�2����T�9X�2W�`-�Y@ߞ�6�'�6�?��GK^9dM�`y��1�6n��~&�§� L(KljjM��JW4��:~.-
����d%�����J�jA�Z����ΑV�l�o̓,9&�HRTR�R�|$�2gF�ܬ�|���^�'�푊{H% P�W���8�)
�"����"�ur臶X�N>oC�1��nl�Ū1��%��`���U�(W/�&�ݯ��Y�І�8Qx��=�X_���yyvY��`9�Fr'F*����C�U�*wk��y39�ߔf��ֶtS�1�@���������[5g[l�V��_�Fc�56	�OJ(���=4sa�]��ϫ�fVРD>�ّr�߁�gO�'9�~y-v?�.���4	M(�[�͍,jxiA�S�
a�Jt�	�����؎~�?}�\:s�Wg���teF���}t���_� ��<ǆ�+�u�ê�P�G����&�Jam|X	f���jW�)C
�=�s<b����
�!Q��g���!>T_�Og���.�ޭ�e	�in<z��@�ƓM�T��0�lO��a��;(� ƶ��a�N�WBDR1Яi���I���.E��{
�d�Վ��mA�����~��0�cVmoT�>�P��ףY!h	}
q�4p���)�H��ʣ-ɭ'O���_�|�f�x���q�q7b�����@�ݓ:rJ�W�m>J���;�^5hٴ�
(`��AF����a�T�p�s!�Y��Y��ΐ|��Z�cfm��l'&!8K�v�Ƭ=�z���ͥx� �W+�1��~p')9o�nN�t΁]>!"D+}<5�g�AxB�e*'gR����X��hWa��^���mX[pQ���'���Y{h���4]Tj��e��l)�^���E�5��B���bU��>��HY}Qe��  0�*����xl��2aLȫ4"��Sp��r�s�����ލ}ٲ=��И�<����xs��UQ܎#8k�~��������#^��]��e��<����M�u$���!��>q�]�zl�LUi���楸M��43��ތ3�ь/�x�'^_��f$���֕�Rw�
Y�9��WhZP������m
�}r8r�Y���7�x����uN.:O|��$l%�����.f'���>m���p����6g�G���,��|�H�E*���U��B^��C�i�����}����
���"+$�.���ښ2�qH�a�ʙ�I���E��DF�%xLe5���� ct��.��K����&bPێ�.����'�ɾ� }!��;�AK�I��"�T��ֵ�q�[�*�:"��yU�:/�-	~~�q�H�\��^=i5-U&����qR`�j�� 7YDʊt�SZ����xzJ�&��
�Ww���;�r,��$��FO�%搻򷍗C?�7��W������Cdʅ�wQ^	A%�`s싐��ؠ���4Nh�i��+��d�m���L�ܩR	���9�{��G@s�����S�ٛ����Шn�xS�(�|
�T�M�������K����P�P;V�_CA�n/
��s�p%�*�����������.�q�C9{,�t���9���v0�ݾ�^XIqR��Ύz�ż�8p7��¤f3��Z?����bv,�ϔ�@/����p����11 �`���p�~�(B�p
��?m�O-7a���T#�REp�JB���\��|���f�_�����y�j%�XF8�0W� L��m"�r�ݠ������'�%�L���^3F@�ᾂ(�0
�K���u[��B�.G�W`P0��v̈́pV2�d3��H+w`[�%�y*q<��w4�Jm�[�v�=�O�X��9���Ƴ����Z^b7��e	��V�'��P<:���;F�q��s�V���	�1�](Bq�
���O>��4�l���#z�(��u~�B�%v����W��>wvd���C��gUm�P��9�ɔ� xQ���x�bfN;Yq4��A#����E��#��Q�W�Kn�tܕKp퍒�TCwm�I��u4�~� ���kdѽ�M3�eNB�sȷ!z.�+{�א~�ߖI�0��F��@��q�7H�^G-������ �dB/qf�?�!�8��K�.��oNҴ�9�f��8�B���pS_�����]J2W� �8�N�@~E�4��� �j�b|����H��eF'��3"��6�\rȻ�$����}+���#R����^�SM���i����`�oc����$ۦ����FvG%��:�
��ov�]��x�[�*���J���On�'��tS�j^O_�{��6�hP�v�*拶=h�>��ɩ~�Hh.h`-�+=	���O[�6��v�m���ŎA���$�]��؃.Ȯ�d+��
$D� d �n�,�yv%w*Lџ���p3�Y�M���V|>Z׉n�.i�cR�])����Ju9i�c@`�󠠢�-��7��D���'����E� b�/w;peP�;eɉL>�@&����HD_w~F-}m�S��]�H�1����3��5���­��W���N8h����.�}��	�5oٴ�+(N�u�����\ځ��M������.�Lr���u�E�A�eb;[^��N��m$��I#��5�<�:K�5Ѥ�0ߺ
�������9P���䀚�K��}O�;�0hݙèGΩ>ߓ�[�ir�Sv�C�e4Nm�f)op�����XD]2g:��o���.O���Yz�6�ݎ!<����[A�떙�)���~�:���u#�x+K�H���+���.�b�:!�-�	fS:�,��F4�`�ֳ�76��c�e;+w
hgC��I�*�����_.&��o�Ε�}��Q�u�����%U���BAerc����=ؓ6���ntwFc��F۬��	^�o��,����8 r����p4�k1l�x"m��#�ك6�S ̗���Ĥ���[��!�����s&���h%��D����2��DvU��#]�J_8jU�h��/)z�_�R���#R���d)̬U�����y��
�S�u^#���9m�9�`�/tK�f
P�9�+ ~�,���0ez,0Y���-�JЏ:QyXL�V���4�b��l�ʛ	��>ِ�O�Y/��jz�����t@�a�+�5Q��E9�˫#�p������}���|��{7�j�W��[�U�Ǣ����x��UӮ����}d��b�݃SiV�ȡ�m�"�U"9����A��Jz1��ZG�����S��e�*�y���a�I�P�&j�����|"L7H�0�b�R^u��Ml��	��k=▚���fU
��:K�J#�G�e�^��n:���O�n�.�E�DK��ߙ ��:(��U�ъ�ٍ�$��%�:_���T3��F��m3���ʫ�c��.Dz]~�f�c����)�i�������ګq���V�x�����1�c�}�|"Ǌ6d������3d%i)�W��K�!M�(���:*���6-��n�����Q�BΔ�4�LK��K�|���@9+h��0#3�}����p{�͘ �g(<�>*m-���`j~�o�VOR<�s:a]��~�V�� ѽ��N��l~;�=�w�R���:��[�����髡�K��8n���t�I�b�!���P����"Dpɯ���;1�1"��9W �Z�%�||Di���C�y�m�MD�v������b�4am�����m4��	!M_!�O5KSwR=FzU��u�V�W*�V��A���1�4�q9Z;x���A����S�U�@Y�s����k1��.�*[,5�/8�1�p/9��j_<��ݯ�gRBy0�*��"7Q�'*J�I!^Ar	jSC ��P��w�I��*4�_�1����\F4�5�{�&B��H�c�7��#v�5Q��=��x3�k��Tư�/�Q�uQS:n�5��ʳ���qF����^�� ĺ�$)dͺ������>z@}+���oݚӨ]������Wh���p���	bx;��q~/?>���H���6p�~�k��gx~�/����s|�[�7/���:����r
U{kjO圑���4	�G"Ht���:	�m�
a���ؐ[j#	Q؃'M�����f��rݐdrX�|�:Pm�5�*�|m�4k��w���Ez������}���C���!.� �
e�"�	���4	��]"j���#�׽æ�o�N_c�[�;��U6��S6U���e��P]	j���s�<�!�F�
�\�����ӳ�]�R���;V1�A?vm9³�Xǿ܋�7dd�ޛ���mg���j���X�w���z���)'=�'�TZ8
	>�k�ث�;�(��]���[����b���I�����Y
Ʃ&aD���R�%�6��(�ϳ��mcx�N4���a�"�h#���#�F�����Vd�7�&�Q0�����P"�f�N-Nù?w0�iKt}U��
���F�Q���Wǲ�!�!(��&�aw��ߟE���ш	Ѥ��B^�E�X��yi{��EF88�翬1���~E�
��������wXAn��fyx7�IH?�8��˹����y1�¶���ʡ�j�n�{1�A����cN��,��y��huۂF�nc�������4�£5�='#9�SO��>�j�i�äE[�k����o��AV���l�������P�Pq;6"����n&.l,�I+Z/���-�}���#'���D^ן�3T^��ł��K��ҟ(���č
GܳntGZ���ۨ�r�2��L����T�E#? ��M���Y�����D�໻�����!W���VG�^:�ٱkmeq>4��u�h� �_��f��҄
�Ք�m�ry�4aΐ�Κ��$u���
��ԩ��u�G�����&��]�����v�T��$��3?A�����Qw�sH�����Z*G�7�<���Z�ׯY����f�&!:�����Cڧ�7��l�S]�HI�*� �F�%a����j:gK|�8y\�1�[@{A�eƨ賤��":�Y�3��JhD��5#�O����y,=� 7H�8N\齉���!����x�c������5�j�K�;�*�a-��A�E�Hbq�u:9?k'4����e-g�t��
V/|Ym�R ��i���|-�bP�Z�����|Ἷ� �5��(�;ju8�訫��4�6I5��4�����ػd�j�$���Ph�f�
0����L����*��,�v[�/R+�9�=,�c�|�%�%�R\hJ���j�'sQt�p����un.�����,��|/h'Ð�]�<�L"�G���!�`�uJv�LF��cJ���|۸�!������5��!&�Ξ�r'����չ�Ot��akЋӧ�~P�~���g��}��w����t���ߺ��ag`��PF����>�m�׃�(�=o��x�Б����N���O�a���'%2�Ag2Y��2��H[jf7��ݦ���7��K(��C��D}��|f�(g~�g��I!g&�gNI;+�XDJ���8����_����ܒ����<w����������	��&$ͣ� Q.����l(M��ԙYE�Wy#�uJv��XR�� }�D[6����V���Ǩ0^L�O3�!	x�v=���gѱ�>P��ۘ���\�\�-CՍ�).�V�|n.���D�h2��2l�Y�:�?�?0�u�e�*�ٮ^g��Uh�}l�K<�Q �Ё�Ѻ��g�PPQz�M�"|Ӌ�k@��]K?�)�����ρ���Q8�N��G��1M߫
ih;���5Íw�6�?&o��u%s����q�6
��gE�<{�.�JZ��Pi��Z����}``3�k@:D)�0r�x��&\�t�y��76�{�(X��z�8_���#����
W��d�m�3���5Y�	"�[6;�#��S��Y��\E;\Oc�-��a	|V��r�S�/�G"#�az�àDQ�R��|��1���"���_c��˺%y���>2�����SL��޲���MS���gpg���vou�^8�G��ѡ<��*`+��t��I�����W��c׆x������HvY���.@+�Nw��6�ڬ�[���~4�Z����; ��:���0�����UKh��x��-�3b+������w����9"ԁ��K�^_t�����*�4����J���8ٴ���D�5���O�Z�'\gh�u��kche�B��-c����>_�tA7�M���)v/c��8z!p�g� ][��?8HP1������Fj���Lx�Pe+��T˵�ر_0,��[��@�XA�>��ȝ7?\��uD��S��jq���̧c/bX�0)�$�.�aE���;uY�f�x�;=�I���t���z>J,ͯ;�ކL�0���i�f�W���!	������Syr(u��d�א�{�yZ~�N��=v�\T r��oH��w��K��	@���-��nD�ӗN7�4dh�1m���A�ݖ�P/���V�9�wOi�L������;�#�tj�)����rEq��'���/+ɲ���}LU��.U[��(���&������1ω�%�}�7�t�b��	5���2��|�+{�i��'y2�p�W�/�n��<���澅9g�����]?g���ٵ��H1>8�8+��hM9'VrK���@�WAm.vλ�KLF��RF'F�-
�~1�'������#}��ah�/�kX����"U��u;�О�e�O�C�����B�nD�yX�*��
�p�AG�G��%}q��d���FS����l�+�|��G�	=����1�,Ч�ږ��?[q���7;iӵvV8��N�/E'�X;r�|/jW�L
\��l[�J��Q!�v��j���A������uAخ�
X3:��e��YkK&@�2:��i$����ynі*7��KS��S�G�9*R�+�z����Qk�<&�q*�q����d���Ny�{Ѳ��#��m/��	��;��|�6N~� ��氩�[N���v�D	$�u�y\a*��Y�l�T\��)�NS��	��q��뿗&~_��}�6���|.�|�3Z`�[��;~��8�_S�'g���;���\�KJՒE3ć��t���f�$?�Sߙ��Ƴ`ʢ�E�:\P+n����f�䡂��c����C���?R}.��]��ډ���f�w�;.`,�\� BI�ZK*�>'���G�&��-��e/g7��Mhw�T�O�W��2��
~Q��C�r��П����w1{�����Y1"?�h�Q{|�����	!x�؀9 t�΂3:��xFo�X���wһ��
��<�!�ŝmm��b�·��\�W��~� �ߛ=��e�9�G鹓& Qz���jE��C���t����/��%F��f'5�,�NR�K�i�u�[hʸ�d�~�U�%g[�~[�õ�B�.�a��Y���*��?�)E��2�r�l0:�vhn���p�Dc��1'�m5�1Ϣ���eDQ�{�q�1Z���%���M�P�� ����Kw���`�m!���t�q�����O0x�|�O�����iFg������?��/�:Zޑ횑3j��2�����42vaȅ�q���Vi%�Ĭl�s�Wk���S�G�&����8���rPr���è���%�H���7�۫����ֈ@g	��c����0ě,����n��ō���淃�5�����w���"yիk9����j&䖗�I�Z)����jdà��[o3J]�pJ�$D<�*�r�H�}Ă���p!�g.+(J%B]���>����9KU���[A�(����oT��?��& ���K�3j���X��YEG�Z�� 6�˚(p:ڠ�g��>g��aB�9�r�%���}�͉m@?� a�˹k0���������D�MOf�2A|��wPt,��p�j8���f��bt�)����>S���5�vQ!���D��� �U�h��q0�fQ|���xh����}���K����\;�� CCuC���_��89sܯ���յ�\(̕D�S�B7��?�o�����l�#�&�nd`�v�3�!:>���7&{�H��ӻ��j��Ś�sS,Vk_=��w�/>�Y��&�Rm'lHm�U���-� E��|B�փWph��^��qN���b�uP6��b����TE_�!��7�g��uL�����@-��y��&��?�ojK{�_�>�����U@�ak�5�rі�5�=\x�΍�x�|
a=`�jĎ�GJ��|0�y�gi�2�d�#�qҮ���ΗC?�M��o`^�<��Nc좶Ǐ��/G_r%[�o�MC�E��w��x����7���*��]_��4;����ɂ*Y�R&�Z�5�J\ac~N�L�o�ϟZ>��R�[���#js��ή0<�?��D֙��]D�;V}��d.�;�ǟZr����i�)�<�;�l[�Gk�k����C�PЭ O��v*�By=�A�a�a���=�K�?�]��ab���Ԓ߹�֑5;zu�Ɖ��K���<�^'n��) 01ǿ���,ΟwO�k�(�<N���T��{n���m�)A6l���ZI���we���BSOΦ�)�`�>�4��sZfGV�[3�OI��jݼ�7IG��
"�d�7wey�Y���I�F�S�U�"�b��L�lQ��m֟Q���AkQ=s^ ��\�5�+)3K8iX�KP�s�\��P�XP$��r�j�?� Zgc?�+�Mj	%s��	��]���A�O%]���i����@���#@^���edy#t���]{?'��|�y�(����߇v%��9�~N�2�"��y���3�t4J�;2��h!+l�Ս�gM�P�%Qp��DZX��U�SH�暒&��%���A�u�&��Y'��s��.��	=` �k~YY^�T��˷+�b�!�^3O2{��?����P�~z��!!/��^,��Q�& "���$t܄����H�M&0(j��;�����C,�k)gr�x˔��iy���0x/3�Z,S����Iu
p*��~\B4�"f;���pS.�����}�$��3��I=���׫��W O!a���C��jFbqU�Y�<�'��D�ʻ<j�v��R�ch�<@ç��Sl?q?ذ��%��K&�b�o��.�d�z��Mӄ)!��@�WD��=2	!9�+}j��GȾ�a�q����5QuR�ǉXJ��Z5�1�B?�ѝN�}��%uA
b�B�Y�~�$�W����NՇ�Λ�Գs?�_tY}�E?��xV��w�,�C_���g��6>�M�at�ح@ӳ���ݶà�i��k��E�\e�v3u��_�.�K�69 l�q)��@��'<��&��y/.o� ��svi"�?1�)mT?"�.�B�D�qb��Dg}B�+�Lr��Y�&�wo]Q�{�e�j�K�s�[�@�z�`�y�.�����apE��_��Q�vk�u/�\/וʥզ��(�����K��� Ć�l�G1T{w����.ۻ��� J `O4�6J]�v�<���s6���d��D��/	FI��R�����h���S�ߞ�����H�T�u�m":�CC����I��gY�L�C��^G��Ft�8f�"� Z�T��6�D!7�����˭DC\_���:!C;�!l?���M��g��q�A����T2/ns�|��.V���x틗����?�&�F�t�9�����)ej�(���}�<-��7�Bx�aU���%��ͿO�=�km'��)y���Ql�z*��5���>�Q��}�]Hs��R�u�S��$��f���� p*Ci���!�z�	��qp/��xW�U���6`j����lC!�]��x�oIf�of��� �眥s�vYK�F�S��/yA���sp�Y������@Ĳ�A�o�<!�)I�I�+|�����=�8ޛ|���h�m�K�Z��j:�쎃*� �w`p��Į�'�U���N�)_�+qV�;&�S��x_����}�1�w������Z*_�W��rj/֯��)9�"���ֲŧ���"�5��{�Oz��<̀�+?�aH��^�Q�d�3.K	�}2l��S6��yP.�3|�R��,^bjMW�KmϢ���1��593DW�6�5t�A���m���8�ފ���u�
j�*��h���f4���b�ۦ��9�̻
��4�;������'��|O3L	l��6��iIL���о��M�c�~�����a[��a�6��ke�Et�����๛$i������ơH������-Q<����-�c�~��;�S���A.��w�s����?�^j�[L9��E*�7/��r#�ܸ1hwr��8��as*y�&Jg` ���U�NM�Q�����n���Ri�)�QC�rxsZR��+H3�ϗ)2����RR8.�F0��/�� ^df���� 5r.�/�[�(�DO�
t��+�(�,L�G��
Ht��H;R4��s�D��cCEUy~�'�S1R�4�߀8/�K��a���H�-� a�E�+�r�N � }��e�����\�F51Rb8�����^���ܟS�$&�ؖ.�6���`�Yh�V�L�e��6r_l�}�0�r��w�GW�{y�gk">J���	|$�(��=6�Y�s�Io!Z�[H��p9�ۀ <��il�eG�w:بi�d�$Y���/��;�j�}:�m�$�6�>by���%�/]���2�uU�4����۾��a�پ���
���|׶�[	��\Q�\t!�H���gBS�P]`͸�����4ߌ@'���z9&f4�����o$N��O�`g)���ݩ�bQC'
�l�-�;}	���?Y���+'0�y�@�pc�Wg�䛡RC7�=�^���rb��c���ܭ1W�z7l(�J��
��#�0����4-6c��}��
�;��g�Df�z��{o��J���'c��J��ٴ��~�%�S'l�]�9���?.-�4r���z��ꎑ�e����Z?~�u��g��&}�Td�int?3o˺v�)��(�{�r���N��Rf�
G�mx�e,����U����uW��b�`��&�/�#Q���#��.Z��gK�s��_>&��J��Zd�$�s�*�ϒ���V��7n�B�aNi�U}&�j��
�S�4{�� p�������.��8M2�N+T�@4�-o��Niv�m�f��c�CtD-"5�����yߵ��ic&0Z�9��� ފLbH`ǁ�����Gj�G͖͛��T㹋q�
����[!~!�V���b/qND���F�6"��(��э�����UYױH�D'�$�}	��C,�Vri�ο�/M0,YE�	Yw�X�,��e���ƥ+��k����S�A�i5O���ՅD-	E`���wx�ITɄ�����31"�\��?w��y>��atd�(3i)��N�0	��z+���Z�s�t '�e�7,�Ǐ�(��L2/�P����Bjk���U	��!t�yce�	�F�"?����v
�kĻU�gQ�Oϧ3�a�����J!�!g�>�1��H��0X����R9Y��M'$���K�*���$��f��AGv~�-�U��Ң;��Z=o=��m���B�?T�^������6!�	��� g��U��-oe�$i(.	P�u�!�!���3�$��ybG��7N�^��n�'�E�l8#��<i4�2��ZK��'Z��8)�9�,�ң�>�Ow�`W���1Wޢ
�Za�K��terhf�y"P���֤}m��2�����-{��!���G�؜�
�PSH���<�mc_�����B@h)��!�nY�!��D��)s�</����#�nPOzK;��f̴����y�m��%F�����̈Y�G��(��t���&�;��������aT
�~( �*VP���!w�Ȁ��!Q��k6敘��0r�i�<Q��D�j���Sۨ�]5ҝG���j�%,w�8,���0�����
�:y�[�L��Pb�aB<�)�U:�r�{�T,C?zO%�R��2�!�K�lt�,�\8����Qx�ek�#�.�}����i���lQ�H�uH��e�co��3�V�Eu��3�E'wR�B(�ί�(6<� ���}M��i�׻c����G�I���K������Ň�m��PP���o�綼r�4�\���Ww+*�2��B��OT�mdJf��r��5����� \���\�h��A��؟�����d��l��Q;g4a )��=������� 5�@	�^i���*f���&C��1#H1y�ʶ�o����^���.�����#����ۮ���+p���gd>��_k���k�!��ů�!�'����t���]�oq�X�B.O���9�����P�^��'�s�h:t��¹�c��1��Wq�N~�%��N�#%�[�ށ��3fXn��Z(����v��B��ǡ��y#_f��ɦ�3%"�@]�'5pY������э�J*�b��Ws�۰���$I?JV#	��]a��.M�� )$9��0��y�����+���o)�Bi�eh��zM
r#������%{	z��p�&�W��w�-ɡrя鍽T���k�0�K�<G��7��Ö&��'0����g���!NO*�������f[m�$þ��y�-Ҡ�[d����W�aS3K&�`�ZW�L�.���u��k��:�.r�7��0,���;�7�0�C�2|��r�F�hz$)r�ۀ�
;6�w��W\��G�Y��%�4r�wOq�b�~/U�D�uf��c~�]N��F�3��:3��_��u�u���Ձ9����������e�@!Ӝ�f�I�ɓ�#���� �k�)��pzEgc7yZ��i?߇y4�dd�)x���a���ku"h�k0W�;ua$�ARz���s̹��;���;g'�ړB5�Ye5�� x"ђ��4��҄��(&��eQ��Y<�~��5�8|BV����B2Dx�)���B"�Hwlvz��2�j7�����uO�H�I�ï2�c	e<w��`xhڋY��������	}�A7@��s��� - ,z+�~m��ҥ�Ё1LpӦAKA�Ʌq�?�G���z�&���l��f����#��/$@Z��E�B|(��(a_�/�z+�x�n��c ���_Y�������['�9S�6q�q�9�݆4���!�� p�ڱ�^����I�����s �E��O��@E��_xGͫ�&b�9Iɦֈ�e�5�ƃi9AK/��Ŗ��K�o��KI��|��2�u�s�Wv`���(���#�h��2���D��H�%�R�h��xޗ�d`5$N�|�q_���-ĭ!,T,��Bu�IJ�w��H����݁�&C�0��l����p���n�r���נ��"��T�0�^7l���$� �"��Ñ��M��NA�4�Q�K1}>�FKiU�k$�[���_��/�x*�w��F��u!+��Ș���:��S���sڢ&�����x�4d��u�nO�c�v7�Z����w�@Y������Eo��8��g����z^�S� �l;x.��1e�ջAL�4Ҳ����s���Qe��o�ab1O����,�:�#:NAn<�k�������Byj����&������{����B��������������a<���x���+F�*��S�${�T��)����=ki ~;A�:���YwD��W{t)�ڐ��8��1@Xeb���vz3t�-��Kh��XgT�7�QH1p�v�)=�2���/�O{���|�U ����,v�eD,U6>(�#��(</_�] D�GL���C1���n���[<$�~�k�o�
~O�oQ��l��˷�Tl%���\��0�.T�*W?�#���a{F��%����r}E����,�l1xW�>I�Ӆ�RWo����_����ʃz�&)���>�v��o�fj	.������W�&�ti˩�_�,{����?�p+��`��3w��!3���u�{�s
�d����[�F5)	��%j����=2t�~��t�l�iu��i#����0Ф9��&�8�p��ylm��*&������� ��/I`�n������?[�$������Ex�б���A�F��EO��/$������j\� ^���P��"QJkI��bq���{��⁀ؙ���ة�E����7J�p��G~�]Q���+W:�
n�����fI��v���������p}�6������L|�䇂��>c����X�D�H|�+Y;_d6��B����g�(҈B/	'
���r�/ۑd�paj���: G�ځ�&>��Ɩ��O}ˏ��t�0A�){=[~t��u�iZ�| �K��2ӡ,�@�nV.�f'�q��e��x.H�Ho�<99ԧ��[2�"��3:+s����J�e~�.A���d��a�Ҹ�K�o5wku�)�7�ӉAl��U ���iUW����&-���%�q�,|��a�E}D�� Nf����җ^)�m��䛱�0PKӮ���l �$�-,� );7�-���,��\�3:��EQ�ms]�� ����asD��U[���ۢ��9�'�A��u�ˏ��Aj7����)V=�}����K�L咛��ڄ������2#�=����/RJ)��]������F�h���]����בX2$���X��F�.�+���v���)�ĉ$�3�J�J�ٷ��}�QPR"�	$/W��I�w
R�E	.HL��|�"�ϡ��j��rww������/'�,�>��k��2��*e��g�!ie�G���#�����'�2C4p��RR�_� OArY
ӓB}y"5�w�@��&x�P��p��bZzj�D��Ć���V=�tzD��ٹL(7���r��\p!hb�
Ot�3�(�����YDajCݢ�߅�VxY�w���Z�e�E���n���c�/ ɽ@���۵$�"���o�ObF�?�)���}���Iկ*^N��\�EW���:���34�Bw��I���w^�r�}�����RFH�r�ϭ
��,�J� ����I��e�S�x�
��d����51���e
㍗{lN*>i�Ll)�'��7�VK�O#�sF{M���%6���K��u�M�Z�7��H���IT���՞��V/ �W;�9C���}Ԅ�A�@\([c����g�֪䞞�>�g�.|�/�i��Z�2�3�.TrV}B�R%]IwR���d	+S	�b��+��m�?H�����
zI#�ܘ+ �%*G�,�7�>�[�|Ys��WU�]�'9U �5��G�lFwj�^�۾ڡ�:���V~s�1���?���P��p����3=N9G7C|)��4= ��x<���m�7���&5V�k8��f����Ӑ�9Q��PnR~;�K�.ȟ�j�>�	Ǿ�u�:�;~�nz�B����m���U��E7M�l�u7�sr�z���#�5�x��,��6�����o���l����$M
��*x>����z!��@/ג!9h.��#�.%�gL�a!Cq.�$�2l��s/�N������8�	��}��fR}�6���Ct���cn-44��K�@}J]�1K�)VaKsJA�0��>YtO��I�t}fSNu�r�԰ݴ=ϖ_���XPmkV�Bz�^������U��w�|��<��Hp�S�������}E�ݶ:����*? �魪=S���xr��nj[�C(�U�Ǻ0�p]�+�������L# fX����5T&T0��h�>��Z�UA�hRO����*:��	���m��'n��ڰ�5�jx�5���a�Y�׾���X"g�u�V�?��%_y�����}�Ny�l�#g��W���唆�<� ��`����ajOk����L���j��@�&dPf�i�!�J��0�ڠ��I�[��!��������1#C~Q��=1c�y	��1�� �u�� �����\�H�C�-h}:��{2�.���C��~W����$��17�.��v���ݣyۑ"�J�YH�z���u��& V���zϡ�`k�X��y�0v�Hl�N��IҀ��FI�S-FXk���%RF%�sl�|n������bd�*(��XR�j�+#�mSd�~ԏ%�C��'���q��S�� �a��C��%��@�`�؁Έ�@�t��i���Ϸ?$;z���\�r��L�%7$�n�� }��tw�'���o5a!=�A����a���Ó�/��jׂS������B&Pƺ�[!�ՍSQ:��~�i�'� B��S.�ę�dR,��2�_��Q�0T͒���=2c�B�K,ۚ��S�[�@-�,�Ӟ���jxW�Co�>�=.j%����&n�aP��"U�}���m����gN��j!<�cP�j��)Y�
�ߢ�G�b!/$F�M��g=@�>�O�������E�Z6 Y�#b���A�x/��F��f�R�Q�Ԍl�r�����8�iq�6񶕲�(��m\��Ԇ�r��8DE_!zlG�N�P����ͮH���K�=��Lf�1�;)�e>	u�ľ���c �"ek�~i@J FJ�
��{���?������ix���lg���9�NVIc�B� E�kR޼��~�����y4�\�­��Z��g��	3�fb�Ðe�&�5t��Q2��2<���<{����̰�^�\x�gn��%����N�v���D"��\{8gZ�*��1�_i4���P2 $�jY��d.��l�j:l���'I�V�Y�^��X�-\(r;?�֒�- э��K�K`�Y�� P
�p�{�>b�!23*�(j	���JK�z��p�-�T����a���Y��Խ�uV���']�b�E�i�܍�j����F�ɝݠ<�6D��pS�4���GE��ۥ*�}����nK�[�$�&�Mbw����?�7��0��P_�2��d�C�s�u�\���0J�4ɂ��2'�I����D��	T|��Rr��I?T����P &�iT���������a����#�Y��W�iry���(���0lC��~���{��Ƀ^������@�l�����H���V�R�H��4��a��D
,y���:ӥ��@n�I(�s���Ow���%�l:�f��"�;�T��5��K�,�jP�7$����3Y�N�����-������gٕ�}�cwG��PR�|�x���5��Gc	�LR��Y���A~����{�A/Ds9n�aטP;E��|R�6����V�6"���^o����)
�V�����̩�a��W��'<��8���jP�	-ņr=Ց\�d�J�'S!E�^:#L���y�����<P\	�k��ot/#��M�l��5D9Y��������\N� ja��TNzq�N��a�ˬ�����X�R��ى������3�tJ���v%�	��@��0-6<���(,{�=�gި�\/�1p:=���G��F� oE�����@����*{��8���2øq3�Z�l���A��?��!��	�L�
�q�
}GK�]��jh�`m(����$�����X���Ъ�� ���<5�����^���-�j�5�	���������L{%l�𤋉n�V8��SI�-_�G�$
	o�����C����<:�i�{9��:(kZ�������e˓������A�΀���ׄ��gx�1�3�
���5�&}��<����g��e�ߧ�������0i�ޖ�mHl:A�p%�-�υ�P��6/Qp��7�2r�b��^�ApT�c�B�{����6N�Q%���E��e�`��5�B��KXl�@2����~!���i1}������@�����#s���,��iV�eZ8woM5n�pe�4֋α��C�e�F@'7�^@_��I1z'�K���%���s�Pc���h���,4���{��6 D����K{�0�iM�p"QۍFN4��7Q5Э/��sVqX�Zt\�����Aڧ�?c��n�+�P��_���L+ʿ��D������w Ϩ)�a�R�����*�_�5i��KI��.�]�W B��r����?�L���G�٤��ع����g��d[p�~]a�;+n��Tm��t�h`C��+�.j�� ^������Ս�� b��&џ�����g0� B����T1��� 8#U�����!3#��h[z�����m�E�u���Y���&� ˬm�\g��$���j4*��yS덈��r�t�kt�������{$����ͽ����
b���[��=
�=�-k��rX;�V��ҵ��.$�"oj`��j-?�(@
����^�w�r��ƻ��v���Ƚ�5:�����ߏ���Y��*U�GPr���aB�r&}/� p�<�K��G�+�������ͮ�Q�@������},�޽��c���b�wܚi�Zy���*�U��b)E�S�r.��r鸵�(�9>*�$��k�������:g���ɓ�nUFN�}�E���ʺHÛ���sz��%�#�{I*̑�7��h��ryv��c��I����b�� �p�߷�k(ܟJ	�*�Ico����Nl;��\��5���_�|O��h|��`������F�7�C�q��P.����"_����	ih$�5
��T��V�\F�%Е���;,Naϐ*�H�����X.Gx |�C��WDA���*H�P.��_�z��': hk�`����ϖ'=L<��@���h�dwv��~��2B�+Sio��"����v�|b����-��5�����u`�6b&u�u��_Cf������kźp���_�xm��$���M{Oͪ)N�o{^"��t[�I�[��!��Y���6ᖏ���fkYS�
\3F�z0,�MCI���N'�e��V#�@ 8Tğsa\[6�)h�xx��1saT�&o�#�su��T�no�j_�����T��)}.��Ds°}kO���FH�m�b�Q��D�\�j��������q��,���05T��Y�%�1�Uni�}zq��K"&=[��M�:2<@�7�۪�5!�_�	B�I��n�����>hn쒈��K�������Rzv��m��;���Z1����sG ED��[����� �"=�df��[�?��#��<���ޚ��|�[9J5�s����3�����	��{��;�i�_�m_��c�#�� ^�qԗO��@�~��$���J!��F0���> T�^y�<�[���=�ϷRR �4n[h\[����5<U�.��B�ͭ&�ţ\34�p-��pF'��Rh��^���ڿ]�s���F}��'<5ϐՑ�3��k�w�����]&Ga���H���^���L�
�SR����y�>(\�LW���{�#z<�U��gV|�(P�����i�1dL4��Ƒ|�Gq>��9���sfߔ?�fD��h���66C/4֬�l���� �q����EՋ��-�p\(<%�n�yc��(qq<Y�hX��t�@�\��$r�.G��RG��sW�&I���Ԝ8.AJ}������[��d�O:'���2�5�����#�A�DC/)���Ȓp6uN��j����Q�4'Υ����7L�b1lrM;'Z��9�E�h��ף���Z�q��3�l������vպ�����ZnϚ���0�f�^����r6�0O��"hl4 M��'�|~�Yq���T嘺�ڮ�NպKg�ZS���ۧ��������T��Z�*��?M���q5P�������7A�>ҳb"S�;�(3�6����ڝ�iU�����#������'����L�+Ƶw�G�����Y�٣����Ȼ���.Ad��/�ѫ ��W>h:��.��b.*t��/������8��Ez�+��q��^�ϼ���`����CS=�%��&`	�\�֟�X��8��E'�mR�{��đIY��&bzJ�%������)�{
���k�h���Đ
�&	�#.�p?�V``\5�V�W�Q��B#'��u����өs�,@��n�C��p�]�nL��@
�pZ<�����+�v���CwX���c�F!��W�(�J�r�l��&�w��UWÆ-���C�Qi��pJ�Ʃ-�u �3����>�퓚�g9��b�0��x�_��3���(f�Ё0x&Sz��i�����r�F�3!G�Q� ��>13����P*�HL�rNy��z9������h�L^�;[�gBO�_F�T%_#rT���iWd[���v�xE���?���En$��Ё�*$lJ)~A�GhM�>8V�oc����E
PI�׫�>܄��Q.���'R݆ )*�=�|&|����:��6�I
�P���]c���9���9A���#Cv�N�׃K�����X�Tq~B+Q�k?ʿ����m7�c�
���kJ�D��c9^����FH����̹����.�>�[�GN��|B�Ϛ�X����[�)%r-y�W���>F 
`24TXg3͞!W%��e��ǃy��hL8���q�x��Ϡ����~�rO]��/��S�/E�#�8�'���X��U=�t�r�{�W������VBk����[�U�q��h�qnU�e/�PqQ}�����tsBڃ��I����R�p[:z�ي��x!P^Ѿ�����oZKI !�v|CĤ*�,�*�n�?�V+)�o��4�7�0��v���l�/z�n�@pk�^��p��}'��%-�[_��q�"Ľ,��A(˼�wtK�|A����P�S`�k����`��Eg.E��K�'S�օ`$4�m���/s�Ҹ�K3�3��*2:��X>F�� �ū�6��KFFXϛЇ��	-x�A�f�tyͥYW9<O*�_o��2ʀ(B15V��7$�d':E����G-Uw����K�PM���Q�7�%@"�)_X��.��g�vä�PN�H�k�i��?�����#�I��{��s�����N�-	�2�7��鐝���m�ѥN�̗�b�;�*T
�Q"��܀��n�'�H4v��Y47x'�3��v�rS�x�lR�pm-g�q��8�3ї@\�\� \�o���?&����޶�0�)M��k��f?r�W~��7:�$��x]�X����%Z���<AE}�n�;��a�j�/i1ۣ�Ym>�,6�le��b��_�k�yiL|�kb�H >	1]�j�����+�c��#�,c��x�,#g�g�1uU�B�`<�W����/� ���Զ�8�7o���	4��g�A�Ϸ�D�,	yp��
G�`��7�Q@��Q:�"=���/>X .�"*���l6nq#����ǻ��0���"�8W|�#�@%��0��/ӡvVJ���T��~\u�\�T�q�Q�(G}�~L��Tgr �݇���x����EĊ�*�;ag?����fc,'�K��V��' {pY�"E�a(3BZ��Z�o	c m0������I��;��ޅE�/��w�u��/vF�E�}g�v����H=��@��m�	�	�l�$۵+Qs������e���\q��cL3�tw�uM�u�t�sͥg���"  1�kR'Ɏſ����wcV A�m3I�ܖr�j�g�n�����J�>Ա�rO��u�+B��Z��$��Q�A=�Ҏ̘����T�u�u�وA���� s�}�ۆ|��=)(�ő#Q��ģ�퐛�����n���'�ҫ�/W[|��8R� $z���*j���n��F)qn���76�nXd(�e��i�ص���׮Pg��y�s�A����%�DT�	�p�Cw�?�G.0�4�;����+�#��d����%�$�}6J�9z�F�|T/�7�z��9߄�jk'�4��S�������4��>�Q-�Ke���e0X��7t̎(���*Xg<kˬR(Ղɤ���0�V�W�Ome%Q3��!:���FΦ7�
:,BQն]oY0�Q���,����O0�N�n�E�PY��B��v5���������^���2�w���O<.�'�ԥ�n>r��A��9����6k��g�r���g�]��E��e��9��+��_�������+F3V��j!H��%fi!nLV�P�`�B��<m�v��u��Yc��mvoيk^U���@�����Ɖ9�*%҈�PJ^�.�(%1�w`4S�< �_����@_f�o��Е���jA��F����U���t�W5#_��� e�r��ުlx�7i<�D�h���lȍ�k�prD����^�)���1Lj�h���:ब�!��X�3��C\��Ӛ`�wZ��s�Х������K͕�F����$�)��,��W�l���l�psԙ(%���*I�W.��&�����s����]ab��d
.a�h�c˪J-a;&��$�%���>��K�����L�X���*	�hj��L_�=�67���}�1�� �_G]���1K�ˆk*|���c�s�=�3`�^#�ôM�V6��Ԡ���0��s4V��+˟���І�x!��vC<��m�7��QK�����r!ʹ��=�l�S^����@W�v��qu��^������[H�{�l�������p�5럸$qg~=[���HS�z��q�w��q��	���q�U� \�+^��A�?�p4d�c�to���6}�ewH��[��E�9{iָ��,��VY4��Z���W��,拏C�_  YH�G\�P�Oݱ�Y�NP&�C4��v}x�m�f@db��'��qԭ��r��y.B����1DK��aB���'U�_��;8Ӟ�|]�����X�?��qDh����Dd�r�:L)���/�dޭ��r�b�^ډ	�*2�Or�K����OBH=�v~}ˎ�U|L�c�q.5�qs��Z��cP��<uL��<�,9f�'��"������Bz�K�p������rC��r�E]*`:v����G�.*w{r���	Z�V4t�`�/
=��S���B�@p|-�r\��.ڦ>IKQۼ��Uԃ��.F�R����ct`�/�%,�پ��̘L�@�&�0��;��Ϫ���I��7�E<T���X�[^*��jX�GߏB�n}:��0$�U�j��s����rCٜ��_�p'�?Cjc�*�FJ�ϱ�Q��q�/!)�J�uz�@B"L���P!��W�p�4�1��v7B��j<fUn��w�ȇ#�j�O�rF�_���5?� :���e�0X߬�-],&�ߡ�u�-�T �&�5նh}��⾤u��`��_X�_�%��+v��6��]b+^�M/'$���Ew�d����H�,:I�L3�s��0�c���O	��%vOް���T���Sb��8]#���/�[&x�ItP�k��[��~F��b�������~����SwA���~-v�/qx�繮|��0ׂk&����O(ܑ|2ci3iU�1�h������n������#�w�Gz���f��Wl��L�Y�MWڑlӮ�>'ܗM������Xn�]��~u?B������j��ďr�1MfXT7��`�����]�}��SM³��E��gh��``-������y��I���-|uqe(��כExh"�0� ����=�7��LP�IŤ���LT+r��ŉ)�[a�Vs�\7:-�����pxxAQv��w��P�n��0 z���Ƥ�r$�0�����\�0���$�vbrQU�`���G�_��J���C����H�ͧ{����ŔI�<�����
��:��5�h���M�ĉ��L��Q��$8�?�^�r�(��y��}�U&e���h�m�|/NɈʵ���[�]U^y���\%[
����б$���5&k�R�~�Ҟ0����z�8����v�U��HF��X�2�J9 �-mqO/{E��وΕ�Y���f`��v$
����܉��x�q�����:�x���� �0�v���z�?Hܵ�A�V����lN����px$�>��\
-�.�[�'}��f�h,f+�N��@����3�=�DzT4p�p� 0��@�T0�Zc�z�JZ����c�G�FU��{�rl����"���Yr.��U;	�~ar����{��_��70NO~H`��xp���p{c�W(�B�]�=��YJ5lf �������Y�f�@B��T�HS�oF�[$fWk2�.��a�F��ћ�ȩ�Ia�%wẍ́����&rZU*_?az�Ε#'aY���A�������z�Ц�7&�ߡ�������=�4Fu{����J*y�b��Dh����\S��"G��e�zǧ�բ�d��f.�͆��)	$I׌FiJ��Z���
H R@e�x��V�R��0$K��ZJ\��_��I��+0�Fqi�,WG {2^�ER���΍
Ys�b�d��7����~�b|��N��w�*F�˟�'!�@a�,[��^�m���[�{� f��R��LYGW~�Ko�MJ�`�:�)H��7��!j�"p\*�h�9ʥ��i�.��F�V����1��5rq���j��D�� �"d�JK.P��%��ȹ�i��R���{ W��q� ���wp$l��/�p�2�gď�����\3Z5k�ȭJ�!B�n 7��W�{�*�.�Bz��ƈ�?�*���f�(���V%�gp1�f��q�<�fM��_zY��h[f�O+>�;>��"�?��jj��۳W,R�]$]��P���_�\�ؐ���G���G�0^�
�K�eE#�vb�^��*�@���#��<\@��}�xP��T�uA)�����*,��,��Q�c��ڽ�a���B�� �������?�p�'v%"��2�4&�-}9$�O21��6�Lh��3���o{d���f�6�>��Jo��f�1�e�ݔ��&�a2̧�	|Á����+{5p��oÉ�Ur����>��ǧ�/��_[`S� G���tD��^�`�d��SoI
0������c��W�ϙ$�����=��/6[ށ�j_�����0O���l b�����5�N␨��k CN�P�ւ�$�p����H�bZ�����Oߛ� }T�j��-е@�p$G�kDC�la�N!��E!�������Ge��\��Oݬ�.0�In�C�'�H���^���@�kg�Q��ϢS��h�3(�w^��A��6�Ω=}S��$"��>��LЁ[��6�qn��kO�w�{�1 z��pVI-�{�(��W��=�Ҿ�~��l�x�P�[,�i��2�
,6�ze�5WWl�Q((����<��q(���pH�ޙ]q�j���4�Ax ���Б�6#PjF[P_`�J�p{m]�+Laxq�t;0P�?W8u�Ln]%�+��-��	N�[g���g��`�������3#⥍�	��5@3ܶ ��+O������1yN��D�$��Yb�<���.�!;��4|��P.Ke���#(5���v�K�^T�k�=eɖ%���Lz)� ^�MiN�se$��ù��+�n D%�p|&9|I���KIվ'���#I/$�=X`���u�L��ʾw28�G���9 i��ۯ����K�ks~$�k��M��j.H���������2�$�����������Ң�dn���#{�WBsȩ���T{��T@���[��Rb�[j��TH+����7�"v�����-���Z�������Sܧ����!<0�|���.%���(��=rs�>�J�������`�,]L�P�VU �3�%� 8X���A"Jʤ��]
��g��8�L���If��R���ɻ�O���sZ���7}����2>�H���٢�t͈�k���&`��+`[=����#��2F�"�23f��T$�hu̵1h�7@dȺr태�`y�>9�g*����xy�t{|0�]UM��#�:^���7;Ͷ�1�Y���$�1�Xy�=O$]�[���F�A�����@�m(̽�s>۵�X7IO÷�Bv�5²]�Dd��Vƚ{	��A�iu���ڽ~,* ���/�����r��J㓄{��(��7��1Ѐ��c]���z�7�����%*H�D��R8$Ғ��G���@����,��>8��<�B�᥆��A�y�iPn�v�l[o�H�Cg����'��Z�\i�S��S��g�S�M�C�T]��|T�B�N�j��пT��mn�[ :5@i�R�����q
���L�c.���9b��J�����C�l�* i2�����=��|h��^��
��<d�;�w��ڛ��6�me��6��i�,�q&0	���I^q��1D��_L���f3��g����ǅ~jĹͬ������A�>,�N|q4>��<S�~����Q��6z�V��z�O�{@I\��Kr+w�� ����y]�A�~N!N�]�fğ`�Ū�
�h��	��A��f�c�F�y��闱��ҴBW	h�åo�8k�go�L��p��$�tp结ou�"�\�1$������XU�^�LȐe������� 2�;_��	u���؍��Љ[ޛ�w�,8o�s��6Њ�&������c��'�9�� xT>�����JqD6��t;� ������������Yv��k��L6�mZ;��E�2���S)�Heˁg��J%r/�ɘ�8;����������n.���j�`�U}��;����)!�LAUK���sop�,0{	�L�����z��
��@���!j_rf���Q0��j|�績���50�V}�!��?^�z�p"ײ����k�=�r�s�FZ�ʘ$ǃ�O�/}o-�}d ��1�n$/n]�sF��Ldqn����#�u�-�0�|DĴu��^��%�De?��>}��@���z'�� ��v� �P1����)5"0�$�[��y�YO}N�^@5��O����>�Ⱥ����;Z�c�ᏄG�oQ�K�|�t�ϻ�r��������%�?����`�\������ܿ��9wo�*Y�̰_�9͒ɥ���;
��l_�Sr A�qO��X����|4�L����ރ�~[�P�v8��¥��@o���V�b����6߂o��M�L�d]��wX8s���{OC$*�؃��C,��'�F���ÑF�� �$����V�=2;�RqAWٚA�o�6���/r����I�{���ִ��@�'��L�Qg&�R���G�2:����d(�V���M�t÷Q{WhL*drZ�|����#��ͽ�_e��D��.Bf,�maZ.ۧ�!�� �9%�D�e+�^e��K�z��U���|@�n'�«'�b^J� !�0�w<���-�x'�B^6S���6�LZdP
ѡ�2�E�	Gԟ���Tq�؀0���C;���PA��9w����D�?�f���*@��6!�{xB��6.�
��'�̫�h�	�1��mnY����3{5B�`�i��>�E�zہ��\�>��i�$¶��3.9������.��"�Ii=�]�m`3h�������{��t�/!�K�*.#A����w��dL ߡ�Y�����U�����C՝se��=���3��;	4��RىY:+.h*����3�2� �l���{��%I�d5�/3�|%x?zU�)���-�!t����f��Sӯ�f���K	��ۿ�����"�C"��6� �oӹ��>끝��;Dp�zM�n�2l�pI��-`4�d $�K�/ w@2*�3Q��$�����,��-�]� <]�Z{����G�����[hG\~J�}�B�s�nW�5:����E��Ml��a�,�\&B���M�״a��%��,/b%2t�놦

	�� �"����C���鋘v�.!��b���O�����鴞�!A�k�.=��n'�/�?�y�A�֥q�*�M����gD�w�%��`���m�9@���q�NL�]�ҍ��-��oKu�Pv�̬�����67l�< ~��}�� ��:spzf�H�m[��o�vl�G���Εj�G��K�|����ّ� #�$_�uČ}����I�ܬwv�k�99�^�Q��}bzr�~���Ԣ�Q��E�n��Ys9�y˓�-�b��OO�9�rRI�Y�F<���*4ߒP@L���:^g�M�&&!|HV�/�RA�� ��[��}�%3�:���{i� ���.BV��z�b�{�����3{i�H�,���f"1�C&�j˂]�g�,���}���\zY���)�bW7T&E������ɟ�X-;}O�(�z�����m�^> �u���J���N�ܓKE=E���~�[�%��h#U��?�[�����?	o\	Y��l@�A��('&�+=����d 0�̏=����F����\��u(�B)�Uӧ��h� ��B�pbV�<�*R��\�ț7�b�������J��q�/!��+�)� �/�'���A.�X%��;�N�=�$R�
I��<셨+���v�ȸ`7Ń��&�SUxPʄ�I�c5�갓�ij����2D��بvA5��S?M�a( @?�"��`�{.�*SO�1$�K!{�!���{WU�Q9�ag݄M~J҈u�Q�������E|��ki�$
����3OۨԵw�	��\ņ`��/ 7Ι��c��O�/P�ҷ���;�_!�⛛Vm�>��/aEQ<Æ&Ӯ��?Nײ��T�]���WW�3�s����ϱn��E֮d��تlev"��gq�.�z���h��H}B�-���t�l?�B�*����:D�2@�L�ɪ]�.XC���"�hڊc,���|���o,��i ,��+�5��FLs��pH=\�|vP�N@m��v��5� '�>*��?+cITC�YT^��R�F.��a�d�����i�x�2���� �M��0�?|���'�qDy��5`{'��%H� o��k�)`��3�/_�+�t�F� �`���f��o�U�9#g�����f��*�ĺ+@1̆�E�����c�2�#L��c(��'���)��x���d���b�iU�0�O0�e�vS ���K��m����ꑸ�� ǔ��bC����Z'S
�B.�����4�MR]��q\��/��8}ː���;��������^x���3�o��z5>@��K���rљ �B���p{8Y@���i���q[�uS� ?��>!�AW\�8jlN��;#��GX���\��k��%�>S�˖�1�ڥ}��U��!S(R���-�Lnٔ�����,&��$3�)��(�Y�;<6��&��5n��}����Ф�]�O'�8>�Ȁ��s����v<n��VkF�P���R��`3�,$�E�r%mcp	Ą
�o&����漌A�l�s��WF˄
�,��i�l��)����X����L��������~��|��z��\hx�UT����92bU��"`�/����c����ƞ� 2���#X4�񖄵ƴMi=�r���o������c�'L�[a�5�0�q(�=o��������٢%�̜�F����b*��&��y��h��/p�%�)�Kj�V�R�R�V2?{�����a��aܴ6V�b����;4 Z(a�JIkK�^�?���~�ne@
���F�o��O=۪���̶�Co���,���yom���ͫ��6� $������IK�Ocke$MHid)G7�h�
$�}�DQ�Pе��G�;G�K�7��ws畫9���LA�0����4�#�h@�_{`���IL�����^��/s��7zK(�z��R�U��ϊ��P�ࡒz佖E��_���O(N�@��_�� �F�����/s/	��z6��ẋk�K�eO�th�&H]X�qc�=��Ӊ{^H��.�ap	R�Q�Y�%�����弞R�T2��㰝��)>4ڜ�E�K/]L(��J�� ��O���tZgm���Ϭ1YP��,���*��9'߁d�u�E�n�j\����P�$�+�;�9��*�Ύ��⧫%�����dj{��X8�`:��SU��$#r����O���h+��7NCk�#k.׃�	���/��ێ��9i�A�АA|�9���jׯр��q�/������f�H |=J��$�к>V��oX%���R�&��h�B�%�8@Yfi�ZQ���\=���T|�'��?�tbN�r0K�g6�R�1zN��6������,j&�����(�����)���0��x걪�G���7�<��Z|by�77�6X|�@j%��%Xz���j��y+�ȸ�z�ÑWΊc�(�3^M��N����S8���5R/����$���<�����^
f�2a�͇����A2��1.����)�]� �d5���QiVv\�(���:�}%��Dq`	�MI2a:e-<��J�7�a}��"��Ēx�_��¢˜p+v\0B���h�0�Au�޶L�
,I�ϦJ7q��^�{t�jHi	�"�V�3�O�'�uu�F��I��
��5V����С�a�oZ���n��(�؉�����d�Q���E�_�������?���RE\��>3%��ܾ
ۖ�������T���|@�����+��m��%<[�" ���ӄ�9��vp��/M��b�L>Q��G=p���n���0ڝI����I�* B>�@7�v��g?
ʿ��h͙�<�q�T"��"1�=e%��޲�%�4�b(�b�Z��	ssVuɺ<�.r��j!^,�Du�Ƒm=>����Y0ֵ�^RY� ��j��:�\��$�_l�2�I�n�	��R�*ǂ,Q艺��'U��<����[�\�(�Ҧ��@�8K�ID�vD�b��Ư���k\; u�@k��wj��c�5��mYw2�!3�>��)z=6��Ϫ��[=q�`��y��`����=��o�ka<���5�UТ�GIc.�߄#�&��uV-���;�����˯��]�f	�Zi�F|�0�k��?�����U�.h��u�����W�״��O��^�3U	.��=1Q���Ѻ�``#I�Y �(��-�Q���P���+@��T�������p�rj���3����*�Hm�����K��9�3+���d�aT��}��n{�5,�G�6�@(���gm��l��B
�,��u-����G��V�����F���M\���k/*�\~#.Կ|���Z<|},��'�I���k�n8=�a7)��G��ZՄ�5��u#��Y�Gc�}�K���i�LG�&�^ЕR�[�ØF�a~j�돜���Zط@�� 2a���x�`{���� �ņ��~�M5��D�*�o���1XG��
�@�;���Rq�ɗ����Nj��<��b߼�T�i������đJ:�Y�,-J�ж!ɠA�{U"rO "d�ⱶ]՞F���}�<�BA��Nn�MѺ�h����b�х�-a'1	�"�L�g3ߟTW�x����C�&{0���b����v�X���D�7�Tf��D�j�~�Z������
�?Yo�eh�c ���X��b�$$���w�����y�2t��"1�)
Ӧ���wL�=��-d�<�	���J���%�m�a�S!�=�%Zp�&)���S�%���}*)jݴ�Gc��k��B�#{2��ŏ����-���K#"�.Jk��\���M�(��RYzB-����Y"��&�#QO�e����!�6xaԵ�s��+�]w��F�3�d`V����p7����Q��f��5oz�'�_�=5��5kq^Y�ӭ�?�ex��m癮m�M���&�zx�x��������5���v��BE�h�,H�����I�8�&������H�h[�&ǂ���q4@E�y8�_�Uxɓ����ly)t�+z�������ڮJ��5VYV�k�@q��V|�	L���C2��� y�����3BY����wb@�߳Ӟ��I �e��Q��
W��� �9�c���e�`�<��Qg.,�.g{N�V>�t�2B���t�6��[���P3��';�JUl`���F�w���/Dk%�B�f�n���3ؑV�'�*]��Zj,�5��_��5K�o2*k��Rk �/f�"E}I\�אL�.d(���㶈`��s�Ko
Vz���
t�x���' �_���O��L�ߍbĺ�@j�	�pb��� �:9ȏi�mn��t�s���n�L����wn�2kBj]�I���l����.̍#|Y.�g�R����TR����Sa�P@oHʋ,�c	7�$�h�f�¢��B�e���W�ن �sx�<��W�EG�/�)J��U�������-��S=��n-;f��?��{�](�5�k~O~�ՙK�ʙ���Lb,��o�h����@z�]t�f[]��ŰU�	�-�d���_����[��Jq<��*����o�,3���%J.V��Z9T�J�ρD��}�5�JZŧ�&Gj���o�5��)6���k�oԥ~m�4�5��܁]t3���T��#
t t;f��d���u&�O�BS�p�S5OH�m�-e�g:г</{Gn.����Xr�~�(��c��C�0�Cr�� �b��	z�5~��L�3�d@��.���Eɬ��"��_���EK�-N����@s'� %�����cndvO��x�9�R��o��脲�c�y���Dx2�}XRZk����U��Q�)��Mk� d��-M!6�e�D�,�����}{/����d!������y�E�4s�d������/��j��;V�E�Bw�~l>uC���>س3�⊤	��Q�J�8�ֱ���y�@Na2��A�ĕ&?S��-���jL:�0�l�Z���x#Z{�K�_0:���D���"����/��}�{���)�D�EG��ֽ:�(xq�*�x�7��T�����N6|0��̟��Cx�(4�m��f�w���-SuA/8��27)�N�Oz�gBϰ�bL�1�q7$��e��� �R'��M�G�(�^Z\3����j�S�i��f��te���*IU|�l����������ӿU�u��-I�5���s���/�r�&ڟ��������Z���V���͹���/�Fb�1-��MQ�}�W�����o�u�:�b�A���>"˵z�]G�?���x��{$�-���DEs�����˵}Z���&m3��E�(([]�g�D���D�^�xQP�ƈ�a�AMk��:���.7��
>��ܮ����4��4N�4��Q�A�K�����mc݋�su���㋚��at̶�Z��k�ǭ�^$��x����}nOn�z��n bZ��W߈z5+Ցd�+>�H�(v-v��$	ɺxV�2��+:�/w��ދ�s@E�$
��+�Pz{C.95Ɍ���gsC�����X�ο+t�/p�K�Vv\�vl�c����Jcԓs��xH��2M�\�}�!�nm�������^)�U�]�W|}�5%��l���! �"�V� >�E/�Ke�zȑ�n�~��Ƙ�,�L��Uyo�<ʹ�耎*�Y�ƅ�VB�.5��o�2�^*
��}�U��9O��1�_��a�{KGn֪���h���&!jr&�b��VS؋��.w���H�T��eҽAi�,^�\��?��+8���-E��+G4��I�@���x��CP��R�ZisO���>{b3�b��.r���mQ�R�a�*�<�D�5�D�O'Tk���*;��v4��&{׋�&���*��p��Ӌ���*r>ؿ6c�(M9"rs��0̈́ܒ��#��x����z�����7�����qE�LH��[<��9�Ѿ`8Uܜ��\>�V�l[�ѣL-��W�����d�'q��z�#�K&��3�\��T~�����E��P��Y��(7���s%eT������
E�F�[�c��W��S�TA`�x�9
C�+5��4���`0>���f�q?�c6 �_�G��9U��x�i������DC�Ot{�J�$�rQ~QFXﺋ{����Bg����뚵bD�Ӯ�@e��<t����ͱݼB�G|����X�0s"�K�E߉�-���Th���8<��X��;��#�IVvβ�w��tM�?���~�PN���9�p� �����vԯ�[�V��_�����X�C\V�l;�x!+�e�AW���/~�N�2Sud�_�=<*�}X����;��Ո(9[i�	A�g8�[m6S���9$�.�1/�g�ncǟ�L/,ɒ��!����p.�k��f�!4�I�B@�2����{a��u�vM���Aa��dT%��躻u���X������@a�J#����h�S%������>l�������OZ%��/�Ss3Bգ*k���ŧ�ZP�F�`+$���x�Zw���@�=E��@�0zO�� ȊB�6?��5&X�zԟK�*Li XGu3L~���ׁȝ�g߃O�+z�'��}��44�����k��0[�b�>e�s\J�ȵφ��")i/��c{S%��l�ZTᒆg��^OФ��':��-R�Vh7核���\|�A`��2t������*�mfV=�]�a'��Uz���e<�Ř3��������	�Lf��C�m!�;gW�?Q��H�jĢʲ�uG��~(rv4�6���U[�5�|�6��je�eݾ���P,���|�����6E{�0����w���b��Q����N���ࣾ��F�x&�#����I/*3��=Ӈؔ����w	է�.�����G@IT�#�h�k�����C�l�w�ꑤ���m0�^VUl��KB %tɳ�纯��9W�����b�%�o'���	���Y�M����qjE��}^�<�?�Q8��~8q���鉡��Ous�v1=�6Ω_L���4�BbZf��f�^�t��&�5�2ߏ�)��P��`=��y����YF�G�$,7��W�Κ[�=���?�G�#gP�r·�y�^6
��"�e��fm�o��%nb�F��ʃ�Ak�b'�e�i�4��](d@��1ݻ�!��:�����@@"=^!ZoMkg��=�DC����.UJ�|vPY^��	�8��͹GE�u�]*� w��K�8D��'���S�aS�w�,qū�8�-Rc�rf���l��J�%���G��jB�Q�K��Q߽L���v?˸��οhэuJ��� ^�n�j�\���8����|����UIf��y%�VK�y�5��k���%!�͇��|Y!t��f��d�'���������i1bw��j&����6N'��{��h����d���D��J��G8�yP��ޒ�8.�����7J.�p;v�� 2;�'�#���3�i�|u=�7�-�1r�Z�giEv�إ/��Q�߄?X��a�"Z�?X\�{1�6xhK�pF��Q���v����5uy�%SJ���4�b���rkJ<o���/��[F)c�GZ#F9�_;t3��h7������]Ԡ'�)�Dh+Z����y %zR���'mۏ\��v�нY�a��I������&T9��ɒRϵwW��"�]�k���ɹ�i�Y	��HG�5iE/͟�\�\�ַk;�����׀%W�y�%C������75�sZ)�u�!k~�X"D||Oi�;��'�}��5����,�>T��<�/^=�m��\4�Da
��`W�'��∨�����"6��#��}�	�Ω���K=�D0_Z�N�?mTc������q�&�>S�Ro�8.�d��'&����_�"���l:�c�Z��_��F�"%1�U. �6-%���ˢ��n��z�QWX�մ�7+���X���%{�#���($j��ؓЋ�ӳ�T����b�oن��`��̶�x	q��J3�MW�f�1'�	�B�5�����ph��QS]f��:��6ׄ�c�yǌH�%�S�)��X�խS�?�w/2�1+���o۰���������J�{���Jv���Kx� ���25���v�P����P0�'�.���I"��`2�O�(%�}ԅ�'hY��_����B�8����-�{��ó�$ۚ�MU{�&$g+�=�8�L����@��]̄�S�h�D��D�� �M�+���8pͻdZ�L�Vn�Zw������������ѥ�k4��F1Q��N�`*�\�N����mgTw�:(\�eX���)`���+�٫�c�g����p�9���2TZ��%��B�������O�B�x��1~���e~i�o�ߋR����]��8�,����Ù���w��}���t�4&�|����5�,9Jr�� �u2o�䁿{)>�̴QUj�b���!�笋 ����].ٶ͂�10�q��
_Re�=����dS�v��w����n�	F9B�n3�����7�)���#��o�ѧ_�)�a�'��z�W���H2}�bd.=Q�x���z�u�Їק[W�6l>W��զ��t�]w�0�W�t��ݩ�z P�[I�(�����(�9�\=_�N>c�	��O����6	l�8�t�)١��ؐ7PM��/v~R��Dɍ����v�+��CJ�`���b\'@��м�})�Z���#[=�x�:��O�3m����fb�5gZ�To,^��E���/`�Q�*�}Gw���Xar�/�#*)uL��h ��w�r�Z�nD���=$��y~4�83��.;X
�����3f��*8X�X�Kښt��7��7᫚���dQ��~k�O�q��n�i �w���#��^ _��u�bZ��T�OY�����P*�kR�m��r��ԛ�0�&�=�:X�\K_e{	=�|����^Qʄ�<��7h�m�l���봁���K�f҉��C��9�`<��qc��L���zȜ�}��4�����m�A�����3X�>�"��Oݳ������Ek�㛄��I���a�*�Z��{5	�1�:��62O�Ro�z%�|�m�N7��I�$p_���ȡ�^7��>X�.��e��޹5�y���#��J�E�r�����"+n�+��d��t��Y�V
�pTXF�C�꫟fb����CarQ��ͻm~m6�����/�vcG�hMB�5�Ai� Ɓ�h�4n��3�}���uuw��L�O0;�S������-����%�o���~�`	�wg�$�w�O���0j�=��	I��+�j4lp�k�L��uJ2��T��,36aG �� q�Q������N��G~9T�(�G �n�;@���Pp0)�z�ה7`/H \�����6Nx���K���$��W�P}:yZ%ee�z�,�����0��D����/"�>et�"fw�g����5)J����}5=���Hu�r��������C���m��}�͌2��S����e�1�J��iK��f��$�"� H�LK��v����@��>�ct��?�X�'~�Y 2ǲ+N��M�/�����Jk��J�DZ\��N�e�����W �5G�U����)��Q�f�3�����z�2s��I��ۘ���V_m���$�c\��L�ːyd�/^��U�i*�|ۄ֞'fO�sqr?�~F���m(,�/|�wS#��]� P���ju6[�������x'��I��D+ł�AO�*�R$ۑ�x��������PW�%��U-�:Ӕ���� .P�˫#��8�Q	���	/ĂK]��^��E:b'Z�Ҏ�D��<���$��v��G��ɴ�c�&Q�Ā����Wp���ְH��0���,��j8��D	���U�&@����ZEZ6��p.�r_)Cg�\ft�#�4����y�������=�#C��dc"ρ�꿄%:�_-a3sD�y_�����0,������#K�&�Y��s�Z�mʓ�U�373���WEk��S߄������_�
�.����Vk��)KZE3ơ���<y\��(�&��a9��Hv3���K`+�zq�B�7Jɜ�!*ЏoϮ�Ys�|�칧/nb@gLs"�!�� �"W����Ogͱ�\�U��N������1�k��ƟCf�޺�#��n��8s��	.Sh��c��ȢH7P��<j���j_��<  P,8�;�֑nE{�qԤ����4�F{���$�ER��'ka���@:Nv�C��d��=��6�3ы�V�ʐ�먍c�9`���B Gk�P9i�&٣�z����;Ax�����<|� �y����4/�����5���f�U������$^�&��yy]�XI�����O�C:���{:��پ���<�@:)�n
s>Z)jc2�#Y��zqA�Q{L�/(5�ZƧf4��s�forn@O����FXv��퓖�\�[h؜W�7r&�Ƣju'H
�8��@�tx<��b�Mi�u+��� ũ+�EB�ѐ��Y��|Erxl�g��3�I��
"������r�g�޴����a��k%��(Bx�m����A���	6��� ԩ�=fz�"�e��.=8V���F���m5H�=�ן3tV"3v���2��*:�cP �p����g��m�~^��tD�@r��Gv������4t�W�s�6��׎)��LB��W�hےi��U&��(��Y{�����X���a�qgtx%��װ�=$~7/3b��4a�ܡը徳�����T�ސt�,�Y��R��S{B��������� ��w��7	���&D�5O{9�k�ah^ޟd*q��S�8'��hh��Q�~�)��	�x�F����	@)*�MN�!�ڳ�����"W���\�D�u��=/Xr.�;�/�n|WD���@ܑ[?!�k�c�zó�h�ns/�@P.����i#�-.���C�d*��߉<��P�d�$�AN�`�6܎Z��t�?E����C��=k�%s�S��)��%,h캳�h3��<pR�j�����a ��U�%�#�0��sn�GIb<6�[�ɻ�d�"�B���{��üKqq�B���7}�U/�Qp���y��Kl<~P;/YY#N�
�A�g��J!�4� O���]��l���"y����띜/����&�/}UF�srlmmKr�P�	p�H�IoS���؞�w:s��w��^�A�������s�*�o��O���5Q!Ӄ|�E
�.��7V:��j9l��^���㙌�"��H,�j�U�V��� � e.3VJM�B�BF�R��^�Q2^+Wd%MB���zZ��6R��ː�&*��]����2�q������%	W�9���,ٗ�.!�%�ƿF�F�=�鿳�hE���6��N@�[��I����y�t3[�0�!~��U��2t���xt߬W�Qa��*	f�\�K�TӒ�a���.�B�
vXxY �A�3�,t=;m�b�ዼ�{��|��.�b\�4�;[��I�m��'`h%�W�-���(d��3��r�i:��ě�
�%.�7����7d��dv."�_�
�gEw/ˊw#��,���?��r�~L�"��
3��<c��U^'�>sTp�OA;�5��:M������H�n}`�t�Lh&c�U��Vb�a�~��{V�mς��+�^��R)1�Y<��pN%�u+�ȱ[��f9ةç��:�: ��^޲�v!��\�h�+K~l#����ד�э�i���*G5Z���S��s�G[�$�m:���&������sgz#�g�6̪8�������d�!�Ò��+�O1I
����Y��#����Y%˺n�^9�{�DY��lv��(K�M�
�'�� ����z�7��m��]��߭U.a�2���+���4FFQ9�"�l�T**��ft��b��~��@\�Б)�* ����	n"w�g�=�.�y�O=L�crP 3�iO���lXL���-�/����]�=uy���M�y��l(;%�)碛{��1��䜫�0�e�7�tԠ��֗��rh���o�2�m��J8J�Jh�{F��;��d�3���g��a��<���	���w��E䦟�SvQ�i1M6c��	M=;�j��Ȟ*�ٹ:aoΙ�ڱf2�0l���|���\���K�o O�F[*��M�Ɲ\!�b�gs�k�$F����*�n�m��_Ia�Z��I'�#���X��p5j	dX� ��y�N@�`��>����K�~p���Ip#���1sR��@yr�����k
!�u�t�;�,��&�1�Dn�ː�-b+-i�,~��i�ɆE@���9��,���9(��n_��5ҟ�X�R<�\T�.T�$|Ň\?���K�B�͸�Ŀ��b˹��/KMo�-�+¼��#g6B�
��6���7c�0�e�!QN0+�t߆#�t	����?TU9��B
��8XF�(�dM�+��3�	|G6+l"��H%~L��УJ���0V����E�X�ߊ`"�s�J��j1��߃����JLcae��Ձ�_�+ABr�S5P����=��r�M_BY?7�$V�U���rW:�^J]I�	+=�J�9n�=+p!de(�_�y�~9y�7�G	��/�*�Pg�R�_��d�bcA�f<���S`��Uc0��V$��i��f���<�0	BQ)-��� �Cz'��sJ�_P��������(�Ul����km+��D�.�P�xQ��+�xh��C1����_�f$nG7y,��>��+�����1ێ�$}o\l������t�s7o���E�ڪc�%|+x)���WܔΜ%)$*-���,��p��e�4y\���+�Q�������BU>�Dm\�>�c����m�����+���I�u��W��z+�A��B�NK�P2:��.C�g��oqU��y���_l ��"�W����}v��@%�a��R��<]G�8G��������J1j7��T.���Ѓ�6d
�8?3�Wa�!��˅�9��A2q��ۊ��~9C�O����Q��i��nZ'��Wq�n^�n��$�[�$���L��.�)�z�������]NK��g=l�~��{J����NX>�o�Q������HGO6�|��"B�W��.�8��Ky��?��ɚMB?�+��e��+g�&����E��ҧ{f���o���먨�>ʫN�̴q��}]Zнn{]�;����JM~|�O�֟����P�/�IRd�����4�/��D��L��c'���|�t�O}�E�(�#�8�,=��n%y�|/:Iig��@�����t����5�ܙ|� ��o7ծ�z����ք��/�t�������dbW��+�����^���^i�/�c\�O���z���ߡ��YʻN�X��Mں9�a�ا�֯V=Y��JijӁ :Q�G��x�!��r��S$l���-Y��>$�0�-�-r��<L|`�pѰKH~(�p$�s:F�(����vYN��uP�� %A�@���{�f[�L�)���Z"*��9F"�e6Ӳ!�V�|W3�{��m0h��C��/E�k����wAip��|��a�aQ��������o���}�O��pz��g�F?A�0Yp|����6;��3�)ywI�y܊��;��{�� n�_�C��؜�t�H���m�������g�{>>��2�H�]G�����[���=���o������H�P;�z祪L��[�Zu��$L�N��}�.�"�Ą�� ����G������~#I�b�C�J-a!&/G-K�i��U�������������֎}������-�v����c���iΐ�d(c��𐷡BPM��9Ӡ�\��6�	�uMYJ��{�+����'��*l�=�'s!�I1�6p��̩�_�T$�r��LQ3�߳y%�Z��š�����7�=����]��l��R���lH=t1��*����k�J��=ͽ���&h+^/HR��5���˱ P����2}H�-_P@w�*b��K08��(�Am��bC��ֻ�F���j_7þi�����k��y]v�4�O�:�3�^g<��O�yū؁��"6;�	��k�n�;bO
�<>��ɜo|3"��������p��XUƀq�q���S�F��rS���@
���+��������BR���m(n�l"��}
N+�F��m[�+v�vg�s)4y�;5�;н�OB6�B�L��2���(-�Z0ԞǴ��"b�u-疦2�5�tɄ1��D{f����φ)��Z`4�����4�Q�e�XUn"��V
�@�#���QZ�iQW�T1,�2N%m��|$x8൓�@.���eX����^B����B�jC��U�l�CX���n�K�����Y�O�����E*��#�Y춏���!�p�h�g��2���d�q1�l�"�����	c��f �:�S�T��
�Ȯ�1�1�����CpVp��S�K�eM�MԄL
X]��cU��T&m�{�a�=�@�Kz���Ғ��wGe�3]75��W�S���w�DPy��f�_Z��f��}�OJ��j}�T��6���m�=4�]{�"d����Ґ}>���j�<Um���ODn"�K]��
X{��cr��GI�rP��X�~b2����E�gN����$��1�Ŕ���m�S<"4��pz�Ř��Q��Q�}�U�%��>p����3�)�R��Գ������#5��ӶE�� �J��Yc^������7
�`����X5[���k��_�J,�L�og2���#r����fT��^ I*ҟ�4  \��
#q-8#7�x(�����H�����}ZQh /�q�#X,��eM�/n�ȹ��ؕ�@�ٲ�Mq�r"�l��h
^��ԹH�K��m�0m,�>����ղKZ1��M���}��ؓt{� ���L8KY�Q�b���g%���Y�{4c�Ѿ��lƾ�s����D�@=�̱@��ئ��9Ok��{��]KC�Ơ�GD��5�G������c�@�M��
���T]ԿZg��j!��bb���箖ddF��Y�1��hFȧ��QEɕPl��Q$��^�gM�⩝�Đ,�z�f(; #��+U����,3�w2!�����>�!�炨C�pt2-���N������#f@W	J���$=OU�Cń�'�{�ꐉv��������Vx�f�8����r#�+�1OgH��;��/�{\���)L~i<���[0��還�:,1;c�uz�D����2�R+QHK����I\���B���$;MQ�'�ܸ��	��U��9�Q���p���� ��nygC���5SI� �%)�ۻ�to��u0	�%z��"��̝�Ӻ�Rs0���A^�˴#8Dߨa*A��4�^�Ԥ���}!�W��ֺ2�psW3���ij0GL,b!�XǄ� �׎qv&�<�j�p=�/��#\�N-��hV�C&d{D����z���cR�0W�Ƀ#]��B�k05]3u&�����/�XDӌ�5�x��B�4AU}0�1QoE��bӽ�~��v���G�K�ǚ���O�]��<���G���<8s����R~��1�f�gg��&���)'n���IC��X���!U�����5��S��lA��6��u��0DL���b@&	#_ݐ8n�����W0YWW3�]�\��u�v��%�;u+���P��<�Dg��?ǳ��#0(�M�y�����签��������&r�}Q��C�Gs��Is0l"�؍��^��rk~���;>D,>�YU���|Q!�]у�^�9��EA�-���_�?�Z�`h�oBο[5���dK����R\I�Ӈ����h�u���)(G�)�1���M��êU�Z�n�4O�B�S�1}�Bf<Vۓ,�!{�C�'��2K�)�����R��I( 3�hE���J:φqƿ���}���醷�`�� �M���Cw�Q�i �{U�83�����,mC����9V�0_4>w�Q�7��a�P�+�-�|�s�(��:ƞ��x�S֪"���F�/\�k������kŸ��gZtHLEV�+�UTߺ���Y��ׅ�ף�+դ���45�1����=z�:��H�r*u�M��4��$���ƨb�ѮW����Bj�����/~Yু�ЬdZ�
�=�6��ս��l�Q=*�A�٠�3�Gp(T��=���������Z��'T� �@j���,����t#�gr.Zv>��*hN$��2n�;VR�6IǛ��Fᝊ�%�='����љ��,lv����ie���P�फ(�d�yz�}nd�� 2�F��6�O�:z�SV]5�ץ敂�$�>�M��e�p�>��г�H��t´��lR+Y�"�6�e�.3�VhXT�P[��=&�e��Z<4���x��F]��{�iF�B� �7�	��,P��ÝՄp& ��l�TIޭ7�]щxv��@�Ҥ�W����xp�1@�|U���s��ǃ�{f��H���a]L�_=
#�T����2�֏�{�� ��c���
K!���ud�X&Z�s�8�AV��y�Xwe�8ر���y����wwI�"�t�9�LF�X�q9Н��L���8z��Hv��Z2�L����4�$���t�;K��R�yN��B�]���-�)J��u���3
/�F!Aw'3�9���`�j�TYST��#�C��0�GY���x_�K�&�Oa&��(��s�@WRH��c�ml rB��W�]#�� Cl(���Yx@�*�$8�W��uʰ��/Z9C�.$������4��Oa27 5;��v#��
(U8X�#�9.�$K�n��%�1�kLP���٘��#�6�\c�O���7���5nb�F�<��UdF�� L��'k8��"k���pf�`��;Z1�kl��� ���=���3�@�&������z�˞^�7�Hi���R�����
�	�����&B
=�s2�-f�'Py���L����1a����Pum͉�6��qf��
�:�-{�ӛ&��;y�Յ���z؎ӹ���� ��oc���G�Ȃ���l&�ŧ��Y��\X/\ٶV�8��H(��ӳ�������YEf��.o�F{�xʁR �q�7,|Z�w�T� ��r��n9��$�_��a;�"�H_�X�� ��,�	v�ӽi~��h
��N�m���ys;`�Cy���a��:P�yQO�i� �EJ�B2;`yEw�5��Ic��(��-�����x˖ͱ�i](k�ߜn'*�N�#��*9�+���f��7J"��Ua>��� ��-,KA�d�h�a|�%��e�>#�e�9WL����bD������t�+xR����������+Nh�!���c�'[��s��b?54M�ɑ��	g&"{lx�jdJ׬��"��*�X.G�#i�Ʈ��xH���+pD��(���؝�e��
"w��L)�fiQS��#���W�C�g?�**���>���5��=
�$�H,��a�}�,kW���������*��JD��TI�?�&!/�!��;�Ї+���o~�[h���`=��J�F�-,A�"�Y����m~9��4h�bBW��י��e����c���!�0G��2�uS����~����F?\���~�C�:-��;�R����G�.E��澺B��4�Ÿ�<�S|M���w�>=5���LO\)�</�W#ɚ��*W���ߧ�J�zF�ǀ��V��^�8�M�0Z��7n�~%��^��>)�7b��i�iKo�6�h�!;�dT �Ӂ����� ���%��VQ�-|l;rq ��
憷��\#v[�$M�tOi�����mt}���ǘ�w���`�|"X����l���b��h;���|��]�t���~xa0�q,Eɮ�TaD��ͨ~h��[�´�� ����-�A�W���.�.��޵�e):�M�E�o�%��FF@5��H��?�븹yi+ȣ���]�#]u"�f��<�i.bT�	�Wt��Vc�L�exCWM���`�ev6�����Z�`��s[+��F潶e�s�y�m�R[r��R�^�n�M*����U����y:�E1{˱�w�<=�8����nl���(�#�ᝲ
�/�0��/F�H��E!��B�|h�,t��"�l�/�����Cne�$�8z��gr���=�`����x r6R��gݜK�s�#���ΥR���meW$A0� ���o4!i��A��Dɢ�>���ᅛ����
q-c�n����2Ww�Pt�Bp̂W3O�RM6��,&(w?�ؕ�U�z�i���"��5��¬xe�3d4�G��f�~��Ʊ�6�=�R4���	{ի-y-��GL��X��Z+1q�����/�����=l������p�'���L��dG>:c�
���#(Ⱥk�qS��F���i]�ߒ�� B��*i��g�`"�&�Po4��|�kO1�kL��7��e,#0.>y���;/�h������0n��,Ic�`)�f��_F,��zZ	WIw����x@hj��gU4V�����������VEd0�פ:���Ɛ
�n�4�rk�uT%�e�'zA5�"�:�h���
�m���C�]؎������?�E�JD��+���7+�¼�Sv�?b�Y�g*��Ot��a���'��_�)�4�=���"���Z1(�h]��Hqn����a��bG-Z��&b�>�r'��n�o��q
:?SJ��KC<ͽ.���WI2?V8�r�zNm��@��,�0��1�����1Eÿ���6�7 ��8���4�B
�T��8H��)c��(b&u%ᴣ ��Q.Bг4�,b�b�PW���ӗbc�p�F�������,ӿ���Z#��L�TVht��vBOŤ�1`@é�����=��]��s�Oq(R8��Cg�r��
w�+��)T��7y�e�����"N�㞞˳�X���J�"O��	��,B�aF�r�G���d��@FV°=ե;6����#�0��^�i��=�8p�͹H�V��xǟ�Æ�}F�����Z-C:�ch-?�»=g�^�'��3�	�Cm���Z���s�s��o�Os+�)N�Q�>Z.�8&Zb&x� NT]��a$R(�9�v��0Y{�C���(�_���K��9���>L�eԏ�M�jC��Pel��K���TG>nF:l�2g�$��?$�Q�m�j���\=���|��J� ��KE�ex09i��6b8�_1/9ߊ�z�J�4�� �~r�8s��&^��Ȭ�I������II���ar>��g�G��o< �,ً�.�`��:��샇sUc<"�m�B�c;�؞^$fb����*�4���_�\J7:��0@D�x�u�\nث����������!��%}���J�翉�S�"\Ϣ�Hb�P\O���&f�a����Z�ϙ�Z��%{�=����j�W^��c$��PF�O_�J-��$	(��ɀ��^b�sݻ���X�8Hd~���X���IF�c.E*�e��CL��}<vԾL5�wѾ����}Gi)���T��E�	k�YT�D���K�K�D�	- �+����_�H��
N/����� K��6�"��;0��n60BV 0Bb.M�珆�&y�����X~�dW��Bf�пf� �O�1����`��ŹK��Ȩ�|5�8�w�����zڛE�nh0�X>� �?h��Eʅ8o�	g.w5�9��М(���f��B"�����n���N�k��&�-s����*������q'(�i��v_�D�)yD�.Pm��M��m��5ʔ��l�v����ТW�ց�OO=y�`�J��"%�С���e3�$���v�$(����|��%��>�A��p���f'S�����o�_H�]T�j��'p]\�B�v�m���e���T\��<���[�k�c����f�q���d}�l��>�]1g���B��UU�ˣ�g:_/
2�#�5���4��,Y�� >��8�"Ƥe�}���oc�7C��f�������":�U�զ�?QZ��Eݰ�DO
B�WV�Lzgc�%�"�R��Lf�=�0S��U���ٹ�>%�7RZ�!��y�B����$�W��u@]}<Di���`j�Y>�n���c4�;���_�g�K�/�8�������v�!-b	�#��(��Q�wz�ŠZ4����>�[g�q
:��o&�������ԟ��j����c��ۛ�-����Ǐ��oRWp�h�&��ԅ��pv��Z��@Ύ��_|������f]P�$@d��`��J�����:V���.q� �Ȃ��U�L�,�ο�K�aF_�V�T}N!�n��U&�z���=�E�St�N:�� ��g�`4��>�t�1�%i�b��i=��.BΎ��� B�i�.�!�Gl]��a�>���I�
:Hfpk�\?�Ԥ�Ȃ
�~�T��?�>2���<ȟ-h)Ln��|��hrS�l=a�����Ng�ﰛ�b�7��g�!}���:M�SJ��Z��U���e�����`�� ���#��c�ѝ����	�vR�B"vY�wI]as<�`0�@�Zޅ�>z/�CiYk+�ה���܈'-���nSb�<�u��$�p����a�p�K6n�X�?����T�q�͢�a@U	t��i:�����Xu�H��ES�	<y\��������b6�Z��o��n���z�64�zIC�(��c�"��p��5�\F�KP(@n�f���q#4�{M�����A��[��=}�
�T&�Ҹ�k�{�q��x�%&�>���*_��d�e�O�Lئ	���@�ٖХC饠
U�׃�nݸU�0��*�[��������!��sx�z�%8r���0���zpz�������ulS����_���r`)*���I�����m��+#W��z�z��"�e�o�=
Y����m{V��jk�]_l���bm��v3M�	� $��w�@ָƱ?%�b��Z�j�)7����X	����UP�/��E����H��\��\�d� ���*L G��
��?�i���)|I˯���*����`7\7�� g"iZ�J#$�:	���c$�_��#�LX��g�H��9��Ь31�̹@�`m�2ς���v�Ri�����f�/��ҏ��eεJϮ��IH�sQ#�8}��-��x�hΙ��rv�°x�)~���X�ҳ�&���E�E�_��v�?�z�O�#��Fiw\�A}b3�q7�:��]d����p�����9���!A?��77BDS��t�	����|R��z}v�����IqY2L|�
��OK�Z,���ۊP8.�& Ld����
�!C~n6t�`���;x��2�@�jܶ���%{ɀ�㔰(�t�gYZ|S��v��!%"5CuR͕|��;�j9��"U��QJ���n ��c���3��Zbb���>�a��w�E�;��������z��ا�gb���۵H��ŋi�M�������=!f&I��<�6��*�9|�p�VxIX_tLDSt����^����7Prs6�d�V����ȻmP�^AJe�^UO�y����W�E}D�$�`��G�R���4���	�/eb��O]JT��̖���������{�b����_Z����!�����[ӎ�b��s-I��Կ*�8v'��_3�w��w#ўzVNIq��Ȅ��@�"��}�eK[I�8�o\"��e��T��W�����"�E�뾄s|#؞�E>gw��d���<y��=b9���M�!�`���k+����{I���	.�{әNfv�Q�*�C�T\ځV)i+��Dn���h,/ok(`���S�ٗmK���2��`�V��j$�m��e<��g�x�h8���T�U�"�Upo�V]��������	ȵ�gw	4�ǣ&������m�^.�WQ�T��q��da��<��ۣ;�>^�뉩��>��]��)Ƣ�`��;M�j�Z[��|����if�2� �YO/�,�.D1v��gnp
i@M�# A|0HBf=���ۦw5�E��(��3U�)�r+Ǿ���-�/ݶf�� yG�b��"׹�h��ڦ6F�W��fE�E���i���&�2}#�nG�LZ���¯g�v��X�J7��tO�ͭ�k�J����5i��q=���{v��?Ƙ�M���"ď��Z�����j1�xG�8"|K�	㛜I2��MG�d��zJ4��2�k�U�yD�P
D��H��7N��Y�q���)���������vA�)C	֛
�ѹ[(b��'/6���`�"ΡT�|�؃�"�B���O�?�C�[�u}�|�1�T+�C��?����5M�i�[����|���(��~���A�;��,ԏ�֣2��$�FP�9TU �=&z���r�R�Iiz(y�L�j�A�f:X(��0��R�C�?欗�$̏@R,@�\�����~�g9�vg�ȳ�/C߯g(ؘ���5�m)��lU�w��*�7a���hNA��T�;�J<w��kB� ���jՕ|/-�D��y�����%a���0"�\��u%OC��q������쯴t�*nJ��j�>RcO�)'��9V	��ź��\1�]�'a�Ci����fP�>���7�}���m싙z��9���w�Ф��� �o���CI�5��}�e9��D7է$S#�.	��^Bࡈ_�K��^��0���s���+3
A�ZV'23��-���-D[��]x,2*�G����˪l"e��W�� ��vM��~(%�)�ڗ`�$4lվ�
̎ƶ�A��c�@�3~�J+P"��H�͢�����m���H�Q==杰�"�*ه��f��q�i��l��u�yR/HX��(��"��	�!d8��7켨���~u��0I(�2K+����`��H��^���JR4k[���޿J�I���+�4�[�{��d����T�w[7�⤍H���O@�?l�,�g�XR������nO�'���8�U�-�fE�>���6=�xuAw��*��<�ܾ>�@w��a{�=���ֻa�P�ShYΏ|k��S@U�:�	b����0%	+̭����)"��;dC0C����<�s�� ��<���!8:¬7L��X~t�j�Q�e�"ҫ�)��w���e����H<S�f`�U�p�2�N-�sz���M}����O
�`1����~ڢ�hz<$�-���\A'�|W�R��Ӥ;�OmdF�Cg���x�am�ߕ�l)�W!S[';
�į;�Cu�~����]�K�q�ǖ@����@ޭ�}�,t���e���*�vu�	)@؝HY�`�`Qt}O�I�W�'�����S^AL��a$���N�|�_-f�81u�?�҆:H"��Mo������6e���#i��Z�OHC�d�+,d��^��6-+��� �y����F���CxM�v�B.\T�p|w%_Y����|��$��i@�f�N��"tb
���ΐ%�Ff+	F��K^_6Pӿ�'է ����5E�p^Jt���S:��l:�m%jV���.�s�����v�¸�ھ������mY��D��7�*�c��D_|"�҇��yv��͏7���9BeI��"V�]��iP���XO���O�f��q��ږ���� �<�W6�Y����gK��������i�k=��n����8���B��^X]�6�q^ -����%@�SM�qJo�Ś�(	MJ���^��(��g#����W?t׹nߔ�^+�}�.�����tԱQqY��ЗP~r�!%��}�p�@���������%"V{"mn��2Y-��Nݑ�̦ثUL���	�s��s�f�������v�z:ORD����i��2��o�sØ�~�t�ː/�i���-ԓ4�hL�p���:�~��qL�X��0����snEt� Ë/���p�K�@v������o���������z&��5*�x[�a4c��v��~gD�8;�X|uS���_�[Sx�n�"��Y�_��DV�����8�#�TS�p�[�=��a_�$��>
Q^�!�@��$d��ڸ4��!"�'�OvP������!���Z��X���l�[���¼���[|�V����"=��/�gp塐Aѩ�Į����4�}rPa�S�]���8ʨh	�Me% ��_�~�����)���Fc����S�<,"zu�r�`%�+�V���zDki��K�I΂d�:F��U�����X'���� �r�)�
�V-.�%ۜa�J�?J(��@Z7�!�MU���E_U�W��A$� ǘ:�^o��L���եJ�	��T O͈�p��/i%H�#{��A:C2d�j's��jJɏp0*��+���*y��k
�$H�3\|�W�&.X�x/\j<tC��5ѨC��F�6NqFn�I��Y��Υ5p��������Nɀ��q{T�p�������g3" E���c�Db��GV���^:o�����lB)ά�H���ϕ��?�MRB��c�i��t{.��s���.\]�ެĉ7q��=��,g}c�A�t�����$Y�Fe���Z��(���Cgr�84s��Ȇسk�dt���:���+B��Z������a���7V�2H^}�}~�\<�<�FpA
a�_~�-�B}k�p_��Ek�#
ĳ|N#k�R�ڝ�ؼ@�%O6�e;�B�j:�unC�Ѷ*	�� ��(~�͎-aeL��e�}\)I�"y0�o�����v���qS�o^�c|E���3�`B�y��4��X�*{��l>��!�o��7|���[��-��m���V:8��!ѿ�ZcB9�ZF!�c�BVG\ڰ+�ԽmE�X�-�U�h`Ek�@A7�|��Ύ���v��T�HL-�o�LjA���oK �:ݙY5�0iR�me,��8g�;C��X����;�?�=�a���eR	�o-9E��\�`o�f�
�\o�!��Ek듭5� �=���S�D�D�� y��Y�6]�,��n6�����E��~��d�q�6h��&@[u�/i�5����� ��1��.?�|S_m�}]�	�!IRA`Wk���{D��]np�r�4cE��*�� |���rN"���	��Q�3ԝawtI}֚w�oM9�g�6#�8/��ި�D���<?�[���Ɗ�7��I�1�T�<E4.�C�Y��Nk��}���̥�/E����蛫��l�U"�ycY�1gɹ�E�y�ź�ΠC;^W��)���%wFn��	e���_�C�]���,�,�n��aAaZ؈��H��� �v�a�uʔ<Zs�$a���Y�Ɔ �L�ѲB����n߾�2�.����3�(�[���o힖��U�����-1<��;�=�z�L^�/���עS�*���s��D|��I6���!������;��щ���:�j���W.e�\�_�	�pᑶתm+��:�����	'�_o���E&�.�MS!�I��,N���N'�e��y̥C�[���
�e@��rr�����O/�"%'2,Q�'��.NĒ灣���uw�5�\�]8/�x�ƿ������ aܡ�����9+y
���z0-jX�%��Kj��4#���$�����#�*��vjs/H��Cz���9���{������PAߤc�J-Uh���,�SS��<�õ�a���|����0�)b#lYm6�>7�Kkurb�x�=�޻�RT"Y�7$���e%h =�o�D7��ϕQj��yɽfDurG��\�ҧS�����ɴ���.������/� ��o����F���e"N|,�Y���C_a�/-�3|��i|.1��{%q�L4m��^x*�`2�W�%X6�
J��}�=��8�djcQ�{����K �I˨"&ӟp��1(�\��H)/+o�&��qG��36�0�M���l]�!o�pyB�j?�:� *�m��֮�"Ӆn±�JJfp%���9f�����^N�Ջ��֊�|������<Z���0K&�麮( ��Y�VGDpb��
��G�Gm(�;�'�(��o������Q﯅,&yE��A�6�.'�ɬ�	�ez�·q�9:F_�+s��nJ�)��I�@γ*G)�H��6{��ٿ,�<g�A��/ۯ�A��K!Щ�	V���>)�&�<����rq�K*l@Y�T 6�֣Ƕ��vq�N���ڳ�IE��V���y���:�]H.�-��
!�'m�m2L|c�X����mF�s.՜>�̸��w�yj����$풘�b"}���i����Xˆ�ҥ(�w9�M���o�y@�����l�Gy(~&|v�l$E&���d5��Ѕ�U!JV�t���Y�鄁�6�i>{[D��~��s[��iZ��0qZ?�8(=ŷ����wg�y��r�K���2dbj;w�[���8��C�y�<:߻�<��#������{�V����,e5��<��yl�R���{K\dM���Z�އB�s�|;X�T�huOV!�[`.^�jS�X
��d� ��M(�n�h}�O|h�h`��WF�6Ck��)�㰺�;�8�/�:�h-6kO��N��(��f�8}T*7��ռkNw��>qU��	��x�/V�[B*��`���\��j�$�Ҁ@w�$�.��H����Y��7���!�/Bnf���6�C*�~�Ӯqn�O��CJ�w���X���I!�zMۦ�����=9G=�� ɹM�i�?0��MM@r/f���ޏ$/܉�~:�+G�n*TKRԀnɖĴ{���[_�Jjb�}���YS�Rچ��ۋU�m�x�#Am���&%����ȑq���<&�7o���
.��X
%���l�NItS܏���X����[��GTK��J��ʊ}���a�>=m�']!��k.���==1�ȏ�
[���!������3v��
�%yT#
Q[?i
u�7�䓻/<�~j�e�!�/8��,�9tFٿU?�[�=צ}�)��9��Χ�����I�ZPY�
�]^K�!�س��`Y��\ �2SZ&u���P���Z��wUx�xOn�?�-$�뜞��R�t�"�'��/��{ o%a�����j���lzo
��(���F�J�b9a�Ho�{A�9g������Y�C��xͭ]�#&�j��6��?��ߖ�i�|RW	��h\xg�d��o�'���$m��
�~M(b�|�˚f��������s�D;��\��n�t�HZ��Mܳ���CB본ek�	����Rz�����t��,��&u�=ֵ��N����Q���*/��g-K����m!k�h���rqm��Z�ïNɴ��h�0���z2��q3�I]U�jV��*^��R6B�й�,��Z[���k��4�	wc�� ���`�34d"�$�Ҩ���kÖ�#\	_����1>���
���x�%6�P�վn!�,x�!H�9S�"=c�jq��0�,��_�x�.�upCq��wd
��"U� ����*ʡ6f;C'wx#F���y����U)��XhC�q����f��ߝܲ�� a{^��>�{��Y�<�s�2#�,C;��}��ʬfn���Z��<>�^�U���s⻐Q���F�O��)��Z��&�(w3tʯ�Y[O�~FAF�����t�n-�-�߳�=�|%~���@�b8sR����$ؑ�z����g�Z�@�lځՍ�»�b��|�@b�oʊ��؇X?�m��mfQA�����VJ/��I��F�mr���,	��=z����dwS�>rQ�&7�%�.�L��ǅ\��/�þ�ْ76�=��q���f�gH�ʣ~��\8��.e��\gcR�.a,Q�a+��	^NيX��,�{�B�+�E�"�A_�h�����4��}���+q��'A�Z|)Ê�O^qa����R�����r\
%���rYZ\�rނ��``y4V�VC�x�"�ӻ����Y.&����u �9e�i�n��]������ �BM[�)�I��{Y�s�B~���A9hz����������=��a�w`n�`Ik�X
D�ZIr�x���@�3/Mu�p�j���&�,5|H��3`�+/C��6	,��b\�PY�� �kNu�j�����]��+AW�@�φ1�~SR���sa���	Y!Q49�ܢ��b�����ѭ"p%$B���zlN!9���~��cu�����˩-�Yy6$\���F6#�|�Qo�<�0��c��H������g=���Ҽ�:�R�Z�E��2s�4��ҥ�&�P7a��IliԈ�u�|�M��T�P��� b�qVq������b��/ xO/o��e���2Ww�����9�����c�+E8���ē`e�n"5�"� ڬp�Tt�i��S�p�v�:�'���5w���k������E�`hW���ѥ+� �-����Bm�i^2q,jw��a���}ot��͈$�eJ|�R�� C��s G��=~�f)R��Y��7�K`IAx�V�B����fq�_��f��O��H>Ueqi�f:v�<&ڑ��:���m���WH��1ުK�_X���ʾ|����yZ��\+E=y5�rM�eS�':vH`��>�৅�y�6�A��cſ��	���F`�����hT�m�����N�D�q��m��w£��R��hu�T�g�f�-��^�Jt�eh[J��@�k�o?oQR�nG)p��@��x�5�-m�(��:خ**��2	���"n�#%?}R�R&�����R�~���.����ǣ;�V�*��4�_�7��������>��U��X�6o��(9/��R�HRU���1ίx���r���m��B��d�F��*Zp��M,���0�/ɽ�Ԙ4V�'C�ɇ(Q7��m�sr���s�H~9:��� 5�8�|�1d�>
�-H�G���=c�Q���3�>�wΪJo�y���Ϭ�6�T��n?g��m��h��d␘�L�G����w��,8���f��c�^%o�Ȼ=j�i]�#�ag�V��p�_A��8�H�7��w�j��1,�^���/=���xjcR���K�Z&e��W�,�5�ʞ�6��V�K�f4;�����,J��W[`l�=L�p���ƃI�R4���L8ϡ�:��~Vߐ�@�q���.i~��,����?�$�k�Ux���)�;o@H2k�G��&{��S/�=��30)��Lf�0�ǍE�g�&r��$pL����z�>�b���p��ւ�rܡ]���	�E�I͐gdzkN��� ���2�r�%��%gIr?��9������+�^�>��ґ:�|��Kfˆ �s�5���BR�{�+w������wfti���&��a�H޴f�!�y"*/��ZL�R:�w���	���e��{��R`z#�8�e�Sڬk��0Gϓ�k��4�8L�FF����jȜ�Ti�9P
m�P:��y$����p"�[�׸��ߞ���F�kB&z�KRD:
$�i�^q9E��~����:��o�J�x@�� [��zP���.�z5������$�"Xy�j��V�O�W�o�����U��4�ͯ�l�o��Q����͜`�3�6�1s� 7��M�[u�~%2���pP^W���V0���;��2��)s�{=�V~���p�j�ɦex0K�lЎ{W�q�\�r`��7~�'y�s��;����t:�xJ~� �����2���,k8o+��~��No��sH8�z�n����:*���'�-�@�C!\�V���������Ei��@�5�9���u��*�>�	�^ �JɳpLv(�"� rOfW�"�01�i-v3�1a�]��X�G�Ð=V��?�a������$�ҀI�^�������ek\��ƌ#M�,��j�}���*!�I�vόR?8�ei֊|"jL�ٷ��x#�]�����!͹m�&&e��JZ��I��k����)	N�%�8
Y��i5H��%Ya����1�N�=l����&y/^^�W�u^�j�{gJ�;��C!��w�)D!�x^�]+R�65�T��z��$#K5#���Q~R�!��9�k�"s6�cB~C�xU�lS�p�dć��(ܛǗ���=�%�^͜3�,�x���9L4a�b>}�u�i�ʪv@�t�����Ȇ_��p�?�+6K>�����M��W�m�Q�j�ٰ}Clp.0I�+�t"H���h�ܚ$@�X\0v�~RZ0.��;AZR�y;�_��>���u^��3V]t�p��s@�����>���G9��:<Ք��ᚋ/a��(�FXO�u�lTJ�ݎu���\�\�-Ի``��k�8�T,_�0^��U�5�Y6x/ܐrO;~5��
���߲���j��)5)��W���l*HnO^0�J���5T
*XB��iƵ��O�\���"�4Y�� V���z=N��4�{0�m�n�	C��~�����Ȋ��mP�qxY��s=��XI�G���Ro�[����ƍ+�Rr+R��ow����"�NC��������<�7����c9�U!�-D� �;W*F�qB��+�k�'Q�|T��|�+a
�[3]~d��b�i�d�?��r��wu���h=�.X�uE�������>��l_��7�36�;�"�.ch�����v͈�3��C�C�հz	m��-T�����A$NǯD[�� ��a��,���E��9S�����nl������i,�%:�NزM�"��u~��1��B�+y$O��eY�F��*�/c��j�������!�D¢��
����lF����\0b����ҽxňUTFb贴Qд���\u�d���!#f��
��e���.` �|@�" 롙6k>@(�L�>q�kCk�f��|F��4����n����)r޳��7�N:�˩"<�CP
��
Sؙ�^�`�-����u�n|mk�8�X��M��bQ���c�Ļ���as�D�%�}4��
'@#Jƾ��Z����	�]��oc���M
���ܿ�}���B�X�7Ӭ���]54�ّجx�"U\�hՆ�H_�Mj7�/�6v���D�õ��`�"�q��+�Ғ-���Ҫr���(�`���E���ǒ�-�B��>�v4���WrԢi�ũ���bۗ��^VY�3=.�'f^Ra0�=�L�΃Z��ڧ�@�Y�#��z��uZ��}#�G��8�\Z�#p2P�T�臷��:�,_�ukl��?&���e�E��e�6�0Ҹt�U����%E4�	YI��p�7dt�iDA��T|B���5YE�7-���L�'�z�o�%vW�v0��!��Ipq�::Z}(
k���k4~��y�6��iJ�Ax����A�}�ϼQC��aAh粴��u裎����=u��|c:�v<DoY���S�9/.c@R+K�*|�y��~ ��@x���N��>���Ҥ>6+@�-�ג���ɫӓ�������RK1�`�!�kۺ�U^B�}��Vw �D�H� ��X�����&�RBG;ri��;�������iL��w ��M��P]�<"O׻r��#�c\�~	���S�҂�e�����#��&�����E���J��4@���=��Vy�S3>�c�0"��ue��I|����q;�]d4�S��Vx�������[���2Q��)c��@>����>���)��u�Р�ߔ�+܊�E�һ*3�9w�,�D�֜.oY,.e���3�h�\w�qzn�r����zZ_�p��$���a�0��"$	 ����}i�G\�ɏ[`�u���q���u�$@̤s�o=��7�>��Lt3	l�f'πYCF�Ş\a�Yo��$'3�Z*Yŋ`��sm�H�!2[��\t�����Cd{'�o���;�ʉk̏F�n+������t�������!X�J��`aү_2{��J��������,}�󧺾,0ɘ�Kf}�Lhj�?����������ſ۸'*�͟�A߅�ϟ���fR%-#2LR�������-bW�>*P~4oe?fy�@�/��TZ�������(4AʒS&@�[8�Uip�^��r������uv�M��˸fg��*lȁ]T�3�:>/q�yU.ʼԥ�N�QۙgϲI9�flH6���Hc�.�#d<?�R�8~:�b�����g�_g��A�wX0S.��j��=��8:HF��*�`�Y)Pn��TO�
&^^rUZ2�2���5J���_x�vi �i�_|}u��~*�����l�.��zS/p��rŠks�rs����7m@"�i뒻��dC� A���`����2kg��v]O8�G\��'?�#M�B/�=º�������gE���ƫڬr�~}�=
0��fϾ��������5O�/�����Dz9s���P��t�s�����!�F@���L2h^�ZW�A��'ps�4�R�2���h��PY��6���d]&+�X:�c�\1y��3��U;�k�ĚGE��n�����-0�l!�[ �����G�a�^M�I�LmH8ծ��a����OtUB�p�ˊB
���F�J��6,�DRf�.��r�}2��Ƌ=��]S��UR�޸^"�0������*�g�{�k:��I�Q�'̽ �z)��ؓ��ϻ�{�b��|;�{f�������1�g�coa�V8��-�ds���So7�Z�*�=~���3;S�E����ΧʉuZ��/F���cI���)y3�Q�D�� 3��+�!,���+䪜@:ܟ��.2��5�O�^�˕��P����7p�c�ae�� ?��I�Q�?ޮ��2�28N�O��� ���/�?�2���`�0�3d�oS�E܅�<��;�1��|m������Z�T��"�o��cr��UpeBt��٠r�Xc���Oøz����X�2����9A����ZG���>�ns�L��D���(FewX;ԣ[f�B�G�L�r̃���/�oQ}�ɾ���x�@�)�ġ�jE$_d�o��Sx̑f�2G%�n\�� J�Ei-��׌[���;�����{���k]�U�7��j��P�.��*25�a�6i�R�y���CM2i���$�L�a�\u��}��cġ�����˶4�%m�Xq��qf�����L6K���}_ӳ�[��1��+�6��1�eyU/:a0�;N{��u[ (1x)�P�j��p��m�N�kց�iۗK0~B������`? #@��ӿx¬C�͈���K�rq����[&Ź���IG[R�Ƀ�D�1/�Sfq��+�L�lo��l=l��#�7%s���n2P�z�P- �32JJ8�Z�p�.��z�j��|{�I����n��J.�L*�R��v3
�22�(��ӯ�2ʭ��H����Yl���~��AL+�`��.8��"���.CϻkH�;�v	ӡ؆����;��bǁh��+N-˴3No���tU$s�|m0)oم�hrr8��5�'ڵ����$Xz�D^���# %8DU_�uw�G}{�Z�^QلW�r����}q�)(,6&�{���T�,�� ~��fF6��(��Tc{��h�%��	�,��m=&_�7��o����\*I˽���Rv���&��9o���=�|�w�l)�`�ȥ[>�t�qQ��βx�&�${~� ��JW�rL��D����S��t;���#TR�i�XI��!v~��AW�}��Z�/n�O������M���#'�6��2	}�FW�z2T�	L�v`rbW{˨��c����,�����+�{M�IG�o-�6��9ţ7M��E��)��7+�)5O�G��]a*`�n���U��6���u\p�� ��]!������)O��J��6�cM$��~�=&�uK��=J�����vƑ��"��:{9���Sk<̬��,٨~<���Q�����'�K��<��u������aH�|�:�*�
~oQci������+�ꨊ���9�}�_�˰�A=b'e�'Zs�1��=|�N�Y(�\��rXF������Q.uˣ���}��RO5n�e"����ǪG�����Ҳ=�>c�~�GGl�%�r��o�w16��h���� c�����j"��M_�^��G-vE�X˖I��O���9���DE~PA�4���h_��XY�fD%�ud=���v��q��Ra�YA��I�
�L1�~���E~Ms��GE�>��~JM�?(�)I3G�,���ֺ|�Q���%�N�.�F�� j^�gm��|�5n:�m,䕄$IAPM�06�k!+W|���m4rI�~3�*8���+���1������f�*3���Xu���6�����6'� ���Kb�$�`[aZ���z��}A��g"L�H�[�z���!��T�N��geu��a�[$�~k.���:F�}�mUq͆����io	k5LZހ����H�W�$�'c���Ǐ���*>\���x����y��Ġ	ö��}If�)+�"�d��6ULs�R�҅@���P c$��b���̦Q� CY��D�齪7P�<��nVJ�č&�`����r���\hG�O+|���cH,�����c8�v�S���9S����m���0�L�Nb�bC�WO�����S��e�+�,�-K�v�4�1t��*��@�L�̯7��A6`(��)�(5���n��T��~c�,�-���^7q��+ F���/N퓠D	AS�kuNr(���OMph�D ��H���(��?H{$!�/�f�E��z
p��ʕibuL���G���D}ML�˓�=1G��?�ȼxt�dh��j
7+��r�ʴ�Y�"Ώs0��l�Jy�����2c�h�g6���o�Mk�
��Ƌ��k��glU�T���t����ƒv��!Á�� ��[V�d:o�\A�vDF�d�J�,'t̫k��8Yo-�������H�`g����B��]�p#T\��v>�P����_��V��Z����2�Y��J�+Z'|	��W�?��n�J۴6��Ψf8'�tDJ��-�0z����+�;K�ƽ�Z��F>8f����s�_� /%:�,�A��_�H4b�7�pI�}%;V.�$�"��K`��$\B����P�r����EA�+x��d:A:}��Z�L��|d��`��1|0�Q����Fߑ�'��,�5��>�ڢ�+W���(���U�T ��Za�6�5J�,�:D��h�/ɚ�Z���
��~�z��)�m��KPw-TXE*�Qu�} �:�\�p��O�{)�������-���@ע��_1�����P�,�b�d�#I�K�H�".�[B�Ɏ�pH�(�D"���j%=ȍHZ�1\o�F��z�����,zs���3�B�d�q��Ծ�V���D��X��Y���`#�+䅌�P#>��&Р��%�F����ZFmp��N�_,�φ�F�9iI-Z��t�ӂ>�;s@�Kn��QۤPkDƃÆ�a�s2X@�����J'�{*P78T��I���?�"��M]|.���Y �7���x��T�S��ٙV7�����B+[�}șѦ
��(;����+_a�@��a��h/�sv��N{5?��חJ�q�d�}�S��x5����8�����^�X� �>����L��4R(���r!�=�r;X��CBrR;��x�c����9u}�0JDl9PL/�8�ÑիhL��mr+��8�-t�۶�gQ��Ŗ+@�Z��<<=�4�)��t��
�[�l���p��f	��)֚,���E�s�x��q���(�_pz�|T�4��ڌ��L�$��*�<£���FEղ����=�p�䒬��=*�f,ee���T�
���H�i������B����z�������۩�C�����B{�t��Pk%;ԥgh$&BC��������v��o�$�: 4��aK֕af�6ȓ|�5�i���c��ͷw�$`H�����;�?<w�b�~����#�N����SI�وC7��G��a!cR���p�s^��#�6HR�Eա�h��o�`K�����#��#�m��'�#�nq��nK[�v�^'��gn{g~�)�f�@
��љ�ɮ���֔��aaΔn�Ő�G	�C6����� Z���oA瞭����S�î4�.S�8v����-�;J�G:>��AO\�;�}���>�hT�,s�~zx�V��FF��|��g�5��X��	�?F�c���a�`|�mL݈~��&��vt/��@��xl�k�l��i��V��P���ZA*����݋7��$�RiG�ΚGqmR[��<�'��/=>�i�����Q�P֓���O��.��[jL\�-�v׊[`d����">_�x�ak\��A�39�C�iv���N]\�<�n���n���^"�Q�I	��.b��'���?<��٨z#@-���y�_y�0�_���%����J��sJ*#��t�|�>����VZ9|��l����4sL]��
e�k��c�Ѩm���øB�T�S�'��ܩ&G�>��&�n�2��l�ѡAo�������:$�=�������G���5�vyʬ��B��2��ڇ_~q��<�X;\%bR�|j$�<n>q�D9}&x)��Q�"�b�7SУB�V�jv�]9��� ���v;�k��wm>ce8���z�Gw̄2B�{�$�xWg�o�>��W���VB0���kxq�=#��v1Mu"�ݢ�C�UD'|iLGP����a�p~�1%�B��6~w����Ab��g�F�� ��=��ڳ�`82��$��o#��s��Ζet�� �K񌭣Ǡz`�ȓ���w� ���{q"��n��E�N�oi_�x�(ٸ��L�]�iI���m�~�����u��fQ�>�OL5,��,6����R���L��ùEO��"Ӵ-�A�p�=/�Aw�(0�$ɏ���/�Tݔ��н���F�	�юͣ��K#ݨIGXy����W�&C��u�0^��eǧ��"��3|PU*͛Y�G�В��z�`Y����� �N��~ʐP��S�qHyK'frz9�����Үe��.J��@�������I���uK�Œ�u��j�������B�?���Xa�~0�iϺ� n�U�-�v�f���=��@X�6{O`����N԰�Y�8��s��۩ۊl�z�n^|�G��,*>^�	�gIz�c��}ǅ<A����mIK�0S���)�,����s��_0(�K��,d�׵�����b�l ��--���è�H{s��Q���J��R#�#�Rݍ�`�#���b�p���@�z��k|"9p��,n�b5�ˆ2U��$bk�b���A�\����ԗ�A|�$;�P�пCR�d]�c��B�X����"�UzL��ՙ��eڃA�5��6Ol�MG�wR������e׳�/�Ds �S�Z5�2E'G
�Z��T+�\�7����p����+*,Ό����^O��R�e�D4P�Wp��-��ۣ��宭y�a�&X��:s�{o�Euv0��	&��_�u��4��gU�2�Mtض e	X��u\d]����!qs�R��L��[�����ñ���j�xߢ����k��As@\�B�ρ�e{�G��q ��2lmVv/~ X��mS��w=%Q�����7���[���1Y?)������1��r��K
|��
g�b֪ؿ��(��O4G�BE+�V���SKY5R�i�Dt�=�2�SB����x�=�,���[���}�A��X.zY���Ԫ��;s����;K��uf���m�gA��\���p<X(�@]6���U��9�>��������
:�'	�׋�7v��f�,r�v%�V�P���ú�N�p���
*M����@����6[)6� �G�v��1�D�<Y@28�ɴ��N2�U�f���J}_LN���i�&g�7�$	�WP�=?�6�����m.�� <�6?%�?��Y���6&��Y0#'"�!}�6E�s_��m�a��g0��
�"}��|����t�W�N@t�-�P�?���ңyC�8��9	H�z�25w�uS�n�$�6Mv���} �	\���${,� ���h�t)�<щsяQ�O���I6�����I̭���!f:�
/٧]��H���[֬�~��a2�c�2�wߗ�v~�D����:�bzf
_�OSB����$�F������I|����G�s�]����������0&�ub캋x�V'a+-)8#�����x�������4�D�	�����.�i��-1�x�<}]f*U�<]"� ��'����N*���'���8�;�(~4To�j\���o6���Q��8���m�sK�����mZ2A��Y��/���(�2��6�}'K��ví ������$A1Fd"�7���v���y������/<��UZuT2��-�� Y�l}�oHR':���B*�8�I^P��j8c�t��R�r%)�7�.f����&���"�E�E���l#�`Y�m��:�J~N_��_��pG����Җ����'H\&���n������޷q��md��pW@�%R(�PG+�0T��X#�o�*�v���~�͡.r�m�2�z˵�A����N���|��t�d/���	S;*P�;`k"y��
<��7�	���������c轠����G�p��|�b�,dG�-�N��z���aA	V�D��*K8�Q�V��FDUuY����9�w�d�a)�kΩY�Ϯ�1S������2�N�JG��qQU0���y��J���W����~bR�X�}E!�d��J0c�?���ᇗ���}�A�1Zh�I�Il6������#t6�G�n�Lʋ�f!;F1���^k5Q��͐�J�>dib\�QsH�S�͔*X�4]�Ns\��95����0���7P�{�S�G�4ݟ\O8�����Im�x���C�I�Qw�Xk����8Y)�X��������GN���|FQѹ��|����"Q�ƥ�����(��ĹǛ��J�S+=��e��YC{�!H��;Yμ�3�I*@;L��WI�qg�*��n��ǝa��Ak�b��CK*�>){h�L�7��Kp�.Z�=F�ݖ�JB��h%`K��-w�m�\��� e����FKzi��^x�c��_���8*�S�T����5)	B ���K��qh�4컖
�2�c �v9�+ �Q�X�yjy�N�_���I������ ���{qe�J����[��X�z2	jװ��A��͐��d0������,'~Cf	H��xT���H`١ ��i@KO=�ʩ�zߛ_.���	��s�-�h�b�_��On�[9z������4+6'3Y{X mO�tf�H/Z��M��Xu2�L%ũ�ϑC�W����"��"����`�lb=4"9�ܿJ,���	��� z���}�r���nK�L�ǽ�"ud���]���]���:�u�\�wK�,�9"n��D~�|����G0eШz���c��cČԊ��O�U�}A�I�WM��!<W]��U����IK�v7�r}��gۃ	�n�O\X��z$�O��݋���y�����s(��Z�
=�g1=�ɸ��K��[̀:EA%si������DY�� ��YS����$���xv>(W`�[$�t�	yQ�����O��\)��XI�Xe�������;����?'�K2�,��*����i�Q����E�"��Q&ЀA�t���4�sMT�<9���'���P�<t99u�܃:#I��/
Wݔ�|뗼�8}��2�r&Ս��5ιۓ�:UeUL.8�ߟ���v:{W�̞b�6SN?h�PE��j���ؒ*'q�~��#%� ���j7UI��]�8����kH���6xh�;Ϧu���Ok�i��FZ���p_H�N�K��6�+�s�� ����_�}Q�G��t��e��3۽�G�=IG�zy��%�/\P�]�X�e�m�_;>C�S����[�g�g���ɚ���j�NN��=����'yX��&+y��	����gማ�� ���JIϛ��\��W���Z��w�RP�����O���ߋ��i��ůE����v���9g��6�Y��ο�;桁�
M�Q�|YMk4�7g-����
�q�DtlR>�anz� ����-�J!x��E\�^�^ �0l=��ޣ�J?Ǆ�z
���-�F���S	z���YG~�ݴ�D7~͚`ߟ�юe]`%R���ߑ�>ޣ� �9��2-��M�cĵB�;"��\�>��v�B��1wH�-��M��)�^P=U�\��%1Ү����� ��5i}�_׿P5�JI��iTqM��	�xXK�b�lz �sfʪEn�'٤��!�D���6�W�X&�K�/E�5-s-���Ų����)�*g"]�hE��#�9�[�y�=�=�.�l��@��fZr�B��u�@�u�Ri�Hi�P#;jJ���J+��W��a�^�G�m`�ڄg?5d�/�J�
]�7�e\��Z�U�����gy;/�J�����԰��Rϥkz�%�2�ᙜKV>V����SZM'4����t�'3��R2�ԅfZ3e�+|���5�|�9�S'c�
����nySa{�1Y�)�u{�?�A��|�)�{�hP�#�k��|Tz�"n��e�3H���	*��ߧ��V㜟��{_l���h����w�5���"V-6�����^C�?���
��&�s�t���e�ƿ-M������o_�`�ڄ-�;�|������E�蟡�W����
��buDAy�[��k��S��Ȫ�,D� &��J�iJ��Ɖr�	�� �ڪEi���9?T+}9���9H{�(����Hp϶���vB���w:��m��c|��q�Õ���`�MM?D���0S���d����.�|��U�Q�.�&��%+`��&�����똌�����9��PW��b�*J�ɒ��GP��Gm`��s�WmO��.=<�B��t9��r+�z�'���O�T}>���㧚+��1�J����GڀB�4��~�]Ȱ]��w[�Y�A.*j!!,B��1���;шQ�DUĊgJqw2G��Q�Z%�H�k$��K4=#��k\+�v"�(�;��dg"���?��6:H��h��RN��!���i�|�5�0�6tqgP����;7�9�����H1L�&�����xT�_VW�TFD��V9S�� ~�/�T�����N�K� ��Gzg��Z�H����E{^����ǖ5���	�^���Wp�/�䣞����Fȶ
u�t
�b=�e(���J��#C�
�Β\��2�{�(�[mL��9��_'�$�٦���MO�FojД�T��ó�0�����+�n�m��V2������ܭN$�m▿?x}���ұ�������>A�Nj94�-�)�	O��������Y+�	��f�R�,�t���w#`�(Vt�y��'Om�g��g@�T3�9��wZ5�������r)�dط��;Ejd����q&�-u/Ǵ����Q<����*�9��i�I�}��H��7`q�,86_=f�yt8aGXh�Q]�&�F��W� {���WHUF�|��̘?������A�v�Gb���1 b�1�zP��QL.�ޟ/���>D�%ݤ>d.�ļ��2����a������d�@����R_�Bud���4NE@λ,ۼ��le����Fd�ep�糭��Hb�
p���o����E\<? ��ª��"�ے	�����_��A�_\am���?�k6u+Yj�u�q��\�A*mN}: �5N�	<�ʵ���:?V7c(��o"��/����e��W-!�:}O�Yo@�sA`&2��t������kQY������hIEf�$œ@�����Xݦ�� ?��:���6�-/�.3�A��3I�?PS xR���:�W�����B��&��a%���
�4�N3^}T�2��n�ݜA�E ��%�,�+,C.Dq�2�0F{k��\�d����k藉>s'7o�ܩX~�=�hD};�A -��i��,H+O�.=���u���Gy���x6�a�.��N�k�F��Ǻ�/��O۶V~��M0�K$n8�T�%%~].>�T[� ��ĩ�����:�F�ޥ�VhT��Ԙ��B�������մL�-���r�QV��%�RJ:D�o$Rb<O�H�������mA���ؓ���`���?���b�����ʆ>Ǻ��9��f������UL(s
����?hp]/�^��}Z��Ke��}����.����|���:�o�Hʹ&�ty�6�(Hz���$��)O��6�K�u�:�@����)ّ�p���7}c���ꎁ�2G��߹��0�a8���ƃ)�����?�֨퓟����ے�_C/E�U��rUwv<�1�4f�4�Jgm�r���~�7�|W����:��8�y�N�O�"���U���x�eJy����%�mY�Gh8"�pE��Gx�Z9Mh�R/���c�3����4��J#��4�]�s�:����U~98�?��n�j���W�2K|���Od���)�P+c��Gn`B�i$H�b됐=�ĳ,l.��?���9h���v����O�M�원����gц�Z��	�TC0zw�G��`�����6z��=��,�$) �ǝ�F%|wΌr/�j��%}{��ӎ�վ/��f�)�˛F��a�PEP|=�����1
Zt(��v�|ج�(IX�{���N�O��Y!=|/�p���D�B!�"K���={�8T��BL��8�[��ѷ��A��R7�"����{�E|�	�V��n��'D�H��wN�x�f�^a Z���C��5��8�F���>�o�?����"@�r)[��\kx�GSDq!�0�@�M�n��XmB����Y!U�.��%(Ηm�n*܃Y��jo�޳C턛���<��RQT؞��ZO�[��VM�N�9mzQ�Q�$9��Kb��n�[#�����VQ9s�Iu.f�S� L�Lc&��/n�U�l��R�٧Ґ��d��Xe<��Ve�@����G� eec�[�t%F��$�s���c�]I�/y�('݋�Η���i��|�o���� 8	ؑ��5�*�;bk��3�ȅ`�|M�2�L��c<9º���YP����'�ua������� o�k\�V���(���߻93��#P��]�PP>ʔ����w�`�̯����Y:�c�*v&lme�d]�.��(�zo�'�9�#��9ީj�,���&<�Kщ�\��%�i��e�|��ZjM��o|�n(/�UO�w�C8�z^�>�J1�$�M�a�+
\�oȰ)��vƳ�qm�At�vw��/�;DC��}����`�+%X<�9���qj�)��b�wH��X�9|s N���B��o�o������Ђz��������~�>yAyRu�p�#w;0q�m,X���Z�@i.?m��@�i�P�lY�,<)�y�_^Q6V��<�2�tb	�ȟ�w��if�v��@�����=C]�����V�L*Ë�/%o�cz���-(@�4m�|��� �'�)��u�f�J�N�y�4�Vȷ�(���iX�mO�+@u'�{\0��
77�N��]�z�d�Ϙ��n����`27�Kn$����U7��kR�0U�~ߊ�iL���T��ߺh�`e�a�������_ʺ���x��6Uh|z���@��<�4��my	����fjϵ�/�����-?� �$�z�]�Pd8�Yi��P��bN�||}pf*K����:�5�[uj��؝��BK����U��׶���D�Q�5%W��k#�!��&�@�����wl��k�]>o��%�:��Ys��C�P��Z��Q`j�kW���G!��(��	wԼl�a�Ye���A�]�O$�}����js��w���+����kM�k9����OT���� h@ί�G��i���Q����}��T��#W� ��������A��[�f(x��En+"~���������r0 ��G>@j�ސF��J���ЇE�T.��8xgZ�|\�����=b��G_�ނ�H�rBISj+����C���a`*R�2��ʶZɴ,�����GP�ժː�A�4,�?�xP�G�/+�V����j(1��uT.Qb���H�i���2�tu��s�`��lV����[ʇ{~W.ԍD�C�:���I�,��ƕ@�0���=i3>L��3	��[�n��_�ɂ
G��RdY���Qq�S��PJ�<�`*�Y�A��r���=^q@�'�ayĉUxd��w�-v�~c�<�4  e-���.a��?E��ԕJq�,P�F�jSjs�����L[�Y�� �����vg;z��������\��S��9�T^��b�Ah���7�q��Y1U:�����XD���;O�!�HGv�q�Ь�����o����B3yPi��_�k����f�4��VH��l�&Ϋ�$��m ^�]�"q���D����+��I��5�JG�(��-���\���r�D#f�u�.�}�����7�-����k��\�f�������LF�t/�d��49��D.'�D���::?}Ňd��nT�0�S_��-�!���'~H�!����R�+;x��l�gq?߃�lG�'-n��8����~GC��7cq��QYɓ�0.7B:5��\E�\�8��z*��� m�9c��	�R�Q�Ҙ/	�V�����۰����X�<㄄��
�������w#�\P�602 �ܑi�n�tn�C�]�WA��S"�\2�x�՗�l����f��w:L�Ƥnԧ��۠��](���p3�?�s���|A�Nn<�����F��ȿ���d�m7���_�s�(�Kes����f���X�g����]1%]�N���ڍy-V�Rm�������*�9^ogM�d��45`�>c}+tG�jl�b~�s���h�nP�:,9��G�6m�荡:%:���	�έ�����$�/���ѱ���G��Hi����Ob[ˣ�Zu�|�W<����P�����DC���u��S/�bm^��/���[̡�
ՙ�O:ܯ�^s1�]v���$�b*>�ګ`Z���Ⱦw�,���^GGb�n�?��vf���p��.���3��Y��1��d�֛M�m�Z����G�����]G�M\�e��#)!Zf~��7>��� #��7��?}��ܗ''�9\{��ږ�e Q0���p��U��re�P�꽪���_�-ф�,� n��i�~��p��	K���@��Yagn�W#�+� �w��6�>�5�~ޛ�����|R3߅2:��;;������<�ً��;$(C;	_��`�!��Ċ���2��k�:њAք�L�p���sQx�e��<#�+�)��$�B=�`R-�'i����w�� �#N�02��DD ʪ��|��O�)�j���o��m)z��m�t
|P�����YR	�%��'�!Z7��֕�ѿ��<Ϡ���%��~/��f��*��}��k<�������#��'�7�Q�9�n�a��/�o�P@S2�nF�o�E�3�.��\��]�S���u���� �|���<�gF��E�:�E��0���.kS���.�=��k(�"�����A�7���P�V���ږ��-� U�%~��Ɉ���;�}�PC*��R�	�	q�w0���x�y�x���)g���y�h�f�B��Sܴv&�����FP�i[q"u��hji�IM��&����&�@�����ꀯM��.x�͛E�Ssf��x�6�}o7}��6�ja@8|!5G���4����4�g��h[�6��A,���	���U^
���v����&$}*%}zt���y(l��H��ad�K��\lN�6Tk��!ҥ}ğ��̐;�V��d����"Q;`~˿)���2ZB(�X�{M^k#	���c ��rLY��wP�e-ǝd��}N�LUnNWNz'��P��j���{;?�f�5�c��j�S�c�gȡ]��v�^$E
�]�^
͎�#�Е���b/���z}^����>����K��Q����8Kj��s�7�3���3�c��vG#tn��,�P;�&�l?v�oog�a�S�t�T����!�q*<[�����	������1�TKyD�S?U��lI�=j�tٲ�˃xh`L vB��DE ɿ㮖��>gz�$����r�	:f�DT����R\��|/�w$����/!\p9�_��(n]ÏN��9���,�8�K7eo�u�.�1R�9�����th�fʊ�{������!wHY�3�U�����}�ĄzG)FIh)#dZ�������~�tX�m46i�"��L&Er1	g�s�O=�\΁������`���<;��ː��U�D3���km� 8�Y;ʲ�cl�2��M/jYm��i�� �=�*6XΥm$>��3%0���L:�K���0�B$�צ�����-��L�>v����8�8��@����:�z�ÈZXo)�+*��K9���Q�g�r��6����0�t��\]F�&F2���]��^� �z봄2���0rc\CC\\��:F���<��U������o���%о�x�j��"��b0u�����ֻ�S7k��j�2{>E�Ccs���cO_I��g�r� �{���%ꗺ9��k�mO �G41���+�ŵΡ�I5;�'᫄����-Z�L9���zT �D�Qÿ��/Z�2D�U2��R2ܝE��[���裌�����x�@�u�>_�����) {mN2Y���R!��Ьe���M�!{��cí��y$h����Y@m��~R��%t���k 
�g/y�
9�e�7�hr�&���JbR�����7��@C�sA��x51<�}?�^,��K�����ei�<�Jwp���<L���F�i��Є0X!\4��U��3{� �\�e�	��_$�T��a���nj,�����f��a�����h����$È*��К��u4A"�VM�U���/�"0��e)����5RT��?e���}f����H&�?8���p�������k�q��k��v���h�o���h�B�1��>F�k)Ya0���Su�Tk�W���6"�N�D���S���D�v ������B��9��Cfz*:��/�Q���:[�0���Ѣ���YMkݮ�������(���B[����8��#���c,I��*���ك�NqN`�(0������m��})����׀�v�	�v*G�����|��������x��.�D�Q�-ق�P��jM��K�h������ݠioR��]H�=��#e���</M<�����=�$�1Xڧ���&�x��]:���x")�Y�Y���-���4� ��<����� ��5�R�<Se�1��mH��v` &$��!�R>�+
���Q(.^u�L�t�����M�v��
�f���Խ��}i�&����Nm����F��z��8�]�ēC͑��bX�3��ʤuV��T���/X���R������X��D��S��z�.��e9F�@� ���i����+���,o\<k��Nc���K���W �RH����h)�Ȏm?�H��<}З��;�V�{H����);I�h�Rʨ�v��TXf1��>����K*X�9�����D��F���J�w����3�6!r�6R(��z�U��	5�C�H���;��i$�K���nMY���[ofï�o��� '4ý3���2���u�����L���f����w��w�w;L,Nĵ�!K@�����S<<�k4q�!~�yH3&����J����̜��Q��H-�M���ç���AǃƱ�8+��j����N`L��05���"-vɃS�}�-!��A���B"z�!~;��Enؒk/U��Hu�i��3B�B ���_Le�uR$O��
���?:��Jr�Y{�������D7ΖlF�@0�'$Qk�N�K�$g�����&b�2Nމ��4���o�7"$l�*�q]���Y�Y�[��g��y��)V?��V�g
,�=V)��D�P�#��:0�o_nC�ʂ��xM��������4���JǫD������ ���G�\���%p�����l�-w��Z�pc�W��,��O�>bM+Z���?4��k�;V [�e���h�MIcw`���Q-��<���T�B���}s����=k���h��໐M�Cr�OC��v
+���><?��,�@��}�>�z��R6��1�2"�ڟ$�@g6��=ZY�T�aN>ZT�$����Q��hdc�j\C��-]He�El�����ن�wG��]�����-ToDǀ@��S�P�����9^�I�ta��m�_��9����!T���1�r�-魳f�
Q���]���e���M��/&	�/d�/�����ӥI���9��K�"80�K8�	�^��ez�!:�g��ǧ�]�3�T�%_��ό�6�s���h��_��箺9ݙ�h;������{��;4�̈7�e��S�ma����G��}��A�̇`TW��Q;��ۣ�����`@_�i����o���C���S���<��ϸ��>1�W)�<�5X�Dh.ƴ��`|�w5F�SL��nC�*�b珴�U�R2�0C~W,7r@ܩf��P���G�S9�n�mj�|7��U�YQEQ"��c����T�MS���L3.��O���Sü��|~Ϧ�@}�����A���2;B}KӴ{��(s�����;�\��&�U�����=�>>㟸B��B�w�/A�,��j��j8��`��ė�61���x�/����b����zx�a�"���r�#�T�JJ�$�=q*ν���#�c)���_�}W���
L����H��;�1d$��h?�Q2�2���mt�(A�Ѝ���~�*�_
��=�������Y�iHMglX�t�'�(/��uԘPs2�E��>w��k^�����*9�	�����T�A��
�d�j9����hM�' � �?��$��&���>��;�mf�f����vӏ_�c�b@2Y��Թ�˾�kj�6�ϗ��=$촻>���K8���^�sf6]*�W9�cG��: j�,�b��{���K��uhn�z���U<��E�g��땗X.�ա{���m�ب��9�O4R�k�*&i��,|%dr�fb�ذ��ݞ���L[�-],8�8S�m��&["�i'�x5,uh�wQj�-�دJ��!�t`o���rvV2�g2/�9��ӟL:� ��E;�>���P�gm�|�|3޴�*��7���֍a�nڱ�7P翺����])4���@����]��C^��r�?�붨�>�7��C:ܜn�6�F��-�e ��6�5�o-S�}�%��`��ll���G]�/D��7&�(��<N ��
�X:�c������C�K�t	�
H�E�A��p:�]J�'�f�[�A� 2�C�n����w��7�W8�X҅�3M|"M�k)t!s��ݲ�1uא)����pl��Y������Ĩ�__p
�_�H��e�!��X�pS��	^1�o�Y�_��	����O�TV�ښ&H"������v.�ːV_ s�>��z��z�%f��v-�9Hե:9E�����(�9���}�U\`����� ����s��iE	�r-li�Q�S��vEo��{��$1RQ<���:�� ���Tp�Q�ta�ΰ�:y��n��������ʊ\ M��Mi6�������4�Q��-���pԶ��Ř�����kB1�0�_-*�]���z!U��z�ɯ��
�>���8���2=x�'�"��VkY7�X
;�epnךݎ���|�@�u�T�{P���SQ���;A�_g.���P$�kýh��Q���6�H����/5�m�z�$L��Lv[Ћp���:?����"�B$��/;h��L��&ZP�%��ϟF�`k΄n�1uP�xL���￟Eo��ju���,�t���|�jU�*�V�o���-�9�'~�"~L s��N'W�C�� ���;���2#�\2pf����[��xڳQt8O��=+фn�/�ѕ2�]�S�,��c^x���,��T����T��#p2��\	��(]��`I�*=�ss«�/9D�,���Z`�X�űB��3�y
���$����%���/�CR�b��*����o�pZ2|[1�W��״���'�=zJ]��~�Y��%�u��ֶ����� ��e'_�!�v�O�x�Jg>I�a��t+�l�jV1z.��������A�<���RA�L�9��?!��<����h	�%qR�FvJ!�/-P"Ϛ�5W/w�aBT��f�=���-Y�K-��JCm�{�ZS<�	�6�<�N��bk��MAí��z�g*�U)�����ᙷ�)��Ј�Z>��X��$;�Hx���[�Q����*�������k�y2 l�� ]a�C�ܟ�U\�ь�M<�ù�9*j[�׎�������&]�+"��۝�(�Jx����#x�7d�)&Q�׈Ux��@� `]u��=V�g����ev����[�}�Q�̎���/��Ze�)�O��{�����D_$x5#�tX��s��D6<�);�����n��u<b�ٽ@PAV�ħ����`Q��X�{�N}�J�Sc2'�=�B!&��#x*1Ue_�?�\�>����cH�������-�r�2��W$����"��ـ%g�cg�����#��_4 ��Щ��t��#��T�>�cZ�4a�����֨�6���_>/�$ щcy|3֝�����v��������YH\'e��r˵�P��o�W�~�1��jROLҸޡfvK�B�nvG��tj��e!C��J+�ض�3_j�uJS9(�}^��S k��d��h�4r��!�o��Ɏ�r��ʘ��������𱫐�Ϳ�J�n	�y;�L�f��~�J��E�
�ץ�ّ�ATnU�-��i�o�J90�T3}�5��n��Ҏ��	z��b̲L��5�pm��*��6��X�)t��"M*�٧<�h�٣�Y�@]�_����Y�eg���0�D����cRA�!�������C$T�w&�����[@�˂;-����Bu��(�m&�y��?yHm�;���\~�SQf�]�a�*r%���6���vǴ��(�����c�8����g�.�W�Y\R�ٮܟ%��)�h9�T4�0��t@Vvp{�����n"c�m#��� �x
�����[�9�>˙mj@���,@YbRΧ��$���J���w���܁�V��� ���piz��}���T�K�bx��I;��@ݪ�~F��{߰���L���#��+G��8<�l�6��?Xa���ӳ�Mb;��ڒk�kf�O{���oP�1E\�$��8���4b&%������]k��8��r;��`�g��
�"�g8tsC%f�*섗Mg.��K�m��J}s�C�Q�|����[x��RP���P�Gh>y ����s�k�{���b�mϛIm`�s;��NB$fnXX=�ӵ~}&RXuj7z�!b���wr��B�y��#��aT'��',�'~��-�aX� ʫC$�R��`	���7��a����.S@n�O����0�`�sa3p���	���%�� TvȗH��@"�����Ne� T���^�\s��~r���b�(Q�!���'F#!1"ô"	'i��QQ^�鍗�WR��¯����̹��]2<5k�Zّأ�R�M���ӳ;������^�'�a~.����Ɲ�����湾H�5�Sڳ��9�)����nm�Cr�ԫ�d���Q�TNu��r㝘,ܦ+�]���M>	�.ϫSZZ���P����[���� &�)�޶�jv�En@(�7�F�{�KZ�8v����ֵ��½]�'�5ި�CC<�q�HDh �6Gs�dX�����y��b��GI@��(�(���V��^��� �t�q��r ���y��²A��Y�J��X�\	7�q�
�Cdp2D���G�a(���(�:���	��xӅF�9��Å�1�]�P�}����m~C���P0/�ʏ`���e>�(-��8�x���q9MR�{����l���Ox��>��у2�\�X�PN`��C$�HD���X|@g���=�ԛ���^�!\�6��@�{�M�ˍ���8�BG�@Ҍ��Y�ADÝ�;����b�]��N6�Q���4�tx�>S��v��6܍0�N
�}�U>t�>�cP�1���Τ;7��JL�ad_�S����s�c�7���=l����a�J��^�Y�D��9E:Kh�҅㾔��~��1n�.S�L�spIt%��|��go�G��C3�6���|�P��uJ�������X<C����BjwaQ
�/�d	xyj�
��o�ok��wz gz���.~6�tF��$�U>84G��!����84|�H��x���^LC�AŝZ?��RK#1���c�冭P�C��&~��]S��N� U�2R���E:B�9��z��"J�UF�+��x����r�Y��Ș���?� HT��-!�#G&$�������ˇd/�,^sD�毦G�F��R�*��X����ǳ���a3�·1�W0�1�F��粑R����`FL]�1H&X\�Em��m4kc�=��5��L��h��@��/YN�v��=��{{����|��}s��<�wut�d��У����fu&N���B�)�Q�Nr����������H�^Qc��`�A�Ԗi&����?u���n�OJ�M	$،�ݠ���kmE\�2�e�A��72��c-�B_r�����0㭷:E���́�#�עt��U۷��UN�uA͞��X�l?I�G��s�~��) +����z���22�w�z7��� Kq	@W���w챝h(p9�dW�5?��j�;��ӓMg��2�{�2�Xz�"ns�(��̙��
"�e㶟o�I�	5�����"H���X�GX�wI�tJǩ��Xߌ���a�ϕN^��{�f����;��I�V�܂ԅ��8|C�̡&"ͽ�)�@)w�]�1�H� v����Nk��j��G5��Z�q�>ژ�ƃ��7_��d�*��/x��&l_�GcR��B������A#�X ^�R�'�L�x�*-�ŷJ;I�w�N'(�`��J���"5����g�K���tT������J���R+N����Bj{h�o��6K^����\
8�dG�E�dn���m����,�Х[ׅ�F�&�Ÿ��lR��nhc%9
��-+p�0}mb����2�� 8U�s\�a�l���q2�����B!��`�z3���֤䇗��8�*B�j���K��>J������I��$MX�mj�-�G��sݼ�b>03Ǻ�kh��]1)��ٺ�B	qU���E*r\�`\=�	�*��ݲ��y����錓,��g]��i���~W�L̍��P�ɝC6���9@��F�i�%�)�ɥY�P�����,�@DA��{L`@�v��ˉ�X�������$Zv}.�1��-��ѝK�����/���Br�7&�u/'e�bΚ�2Ȫ�
�#�27N�q�⺇d袞m���Mx1�6r��`��ߺ9�!�sH��<���+����Eqmq�5�u�7�3K���on��b�6�kY��̹���$Q�>/Q>���u�pk��e��j����[�,�܉��SDY�p�N�B�7�=���c��ˣ�G��[�q���l��l�^cze�Y�Xw.��B䴧G�`��
��.�P5�h�
�# �I9m�c���̸#)w�����࣒�!���YN +�8X;Z�O�C���IO����v�/�+�Ϥma:�˅d!��D+��O��F(���XO�%ͱ�,~M"�2�O|��8W"���/k�g�]}<"vWn����Ds�Oc:��L'��q��[s\�$��Sq
�e]�s�v����:�\�Ў�o����.d5o�̷��0�v�Ss�ۢ���p���+��x���u�p ҰFϪ����-��H���	��C�:`Z�n; 6�'z>�FA����)�Fd��v^�SɌ����s�����K�#\v$�HH`�z�X��S5J��Q����p����w��-l?��6؋/O��K�����p,7�K&�F��*1��c=|��7���5�MCJ���n����:50�Qs�:A(PO�q7��Y�/U.q8sa���m�3�:7��!`P\&�s6�B`% � &�IiARt�Ovl��W�8�P�V
pZݯ�|Q��k&��&��~%�g����Ҍ��fm���HPш���hK���*p<�+g{vS��ɟ]��+�Z*mP���fM��zI�@#.Hq
n�d$�� �u��ٕfpx�?`f����8�?l���j0��o���RT�x�����n���̆gY�-�BBSK���Orn�āU0�*�̇,�eC�4t����F�Ed�e��U��%������[5�]#r~��A411��1��:>�cLSn��	;�'�>ۙI�9�~�����ޯ�_�����v
��?Ԣ~�*>��u3�NӗN�p�ƣؙaIy�A�no)£V	R�a�#J�#�:�ʟ�F�MB�a��zQ�#�խ�%%"}���ןf	�LjȤW1��+W�?|��NOO�
�ol�T�����%�8k�����s�9�ߧMY��99��lԵ�#��)��~2%y#�%bhWB37�L�Q	���/ɺP_��{�@����	J=��0Wx���G<}u|��Z�f�>P�y]�؏MbA$�VVo|��60�0\���\�>z��f#��M����손c�#@�H�W�#�ܘʷ�oa�0^�@�������b��F�ra9�g�)�)��ϧ���U��)�)�]*�#vBg!�$r�V�ʜ���q����M��X�7�]�M��F���"W��K���o�G_��ɗƲp�� ��B���5��s�m��B�B�L�%���C�:��v�����q��_%a_u�t9%W�\A�U���z�C�����<��A�z�p��a�{5GMVLK����x,R�G|K<��XY��%8��P'X���/�+�0n�F\�$�H�Uݐ�P��W�æMN0F��O~��\����,�����W����wɖ������Ͱ������"�Xg���~�W���.����������^S>�a$5k��`��������n�id}�s�I�A"SAVc>��!�G�M���J�i�E���#c�������3?z��:�  �Q�7�l���
����{z��zG��
Qh�]6����s$4�aBWo��x*��Tf��[>>�ڟ�O�XY]:��q�D��Q&=���T�J����՗�N%D5�!ǖ�O������Pix "��	�+;� ��\����>��;�\�'�6��U^��l???,�(^A�]��0^6C�"���:F]Ӿ{>ZsO�W�Q`z�b�m�sd��壨{�{�Ϛ�\kƁ����wȗAZ�ޗV�rBhfwq,��]i�c%�N>D�qfd0�V��N1j�TNa�H�3j�k��k):����y�2��'&�n�^ɰ���1h_]m�E����Ea�c6�#�E(��)Xv_⧅��M8?��h|ح���
�tU�x�?#����=���f��$i�8�H�qDkMᝥ�;<9)E�6e(�O���\&<S�H�����
|��9~U�p���uD����sL�F���q�ޞ�
7�P���q�@�&�*�Rg��^pL�b]�9������v�EMg9��L���(��լq�i����
�{��o�����������P|�#�+��$��Q6 � �[�7<���,mP��A��Wޚ���
, Y	_�utU��9�w��6�/�<B�pZb��֮����5m��iE|vvF��*jhɖ4�x6h�3[!ƛ&>��q2w�.�*�W"K�X��7��]��� �O���Y�O���x�~D9�D���c�������c�L2E���/]�Um�x!̧W������@O�F���7Nr=����ڷ,K�����B��j�i^>E�������F���o�z6���q6��@�HA&>d�����g�1l1(�3g����(�<|_��"�ƿ��M�Y�T�]>�7T��}X�.K��H*�S�k+�2i^$���������۷��Q[ ����ue�ӕe�z%<-Љ�b���.C�Tb�G��g����xy�����S ���5�$Ee}C�)tQ�ա��.t:0/�t�PB0���������8J�#��C�3>9����ͩ�ƃgҾ�t�m�ˌ��F�ڕZ�U ���>����X[t�@�#4��t#��'e] z�X Œ�(���f��s��k3=�M�H�(O�G�t+E�������E宇 �R��}�<�r*-$jp#Й�XcamTd�ch0��C�L)�f�H�z��e69�(���q0���W�������R�6�_�Sk�g�k����P��Y�I��d�5�W�����@���� ~9v�څ��X����?62İ��j\�&�h���ћx�4̀�d�|d���W$j����6�]�V���������6h��O�����S�3#M�'�ڇ&,4ϴ�
���W����.���y��K�Y��$�g%W���Há�J�sǼ�u�����H���e���/���r��ݬ��ѽ|��Ǐb9X+�A�⪍�͖�և`2�`~
�",�We��wj���6C�y@���w�.}��7��ZU��w�QtLƭ׉�(MKG�(��m�҂e�36!�e�ܼ�W&��J�!�$رʍ0n���W��	���[s����:��C�Ĉ]8	k��J���*k@�n��!�G�& !1Ȉ�U�BD�J��f�k^�lW�f�%�W-��t>q�F�E��g��*�
�F��1i��&��nj���6�I�S�.Ta�Ko%�j�fu�ɕW��G�^�P��%7��xc��X*���z��	�Q�ZR}g��@�^�2�`	��P�	k��Y|Q�o���%>!Yl�����2�a������A{L���ҭ�L%�
�鱠�!��"� }w��t���0[\�鏦�]*7��)(d�F��Fy�~r!7l.�v�_B�+6�����"��oT4U���|?	nɴp����
��(��]�u�,)��΍��{�c��n�����>K%)f��uP��Ty*r~�c�/� ^��h�pLq����$��׼6.)X#* M�3f�/-��7I�1��$So�X����$
��S_M�/{��= 1?��][�Yֶt7I%q��0�!��*P�@�����Y&$�D�?���NU�^]�R���s�c7ƒXN[(jˬ.� ���V,�>D�!I�O��q����Cyku�4^���a0����]�N���qҞˌ����΂9fJ&^6Wft�
�32�ʲ��b�g����䴃�Ԫ���܏����Դ���'�9���S%�ӽ���>𫓒�^��aA2�)9q'�)5˿X���DKc��E	�L&��[��1��L���`�k�T{��9f��ퟗt�����@�Ml������̊� �s�bH�?|b,��kT����;�KR�#�m���?�O9�,]��/F�,����N��B���|Q���܈z�_9��ץ/�ȕ(9fķ"l�|�{Lw5w�W����&(��9�>��#�MI;��lP^H/�G�Y�t-w�*<�{�c��j�g3��@X��5S�i�i�
���}?Ƙ|B0��k|�1ϣɚ5�R��Dj�}_��'�����9�8�pIr64,�8�O�FK��cj(4ªx�t�Z-Y��b@��f߲^̃qi'S�C Iz�K���}@�u1��{���"�[_�z"}�����Y�b(���AVH��TY;���_��FCFȇ18z��l��DAP�1�+��l*�T��h�����U���%3���	�f�d\{�"�s�ԕ��M�%���s�\J�A��/����e��i;Y�x#��O��8_������,��#R9.�?ښ#j*́(��������^%+H�r��	{@�c���|�j�/�q�Ln�����5�V����Ã�q�Dv�C�����As��R6_��z�yd��
8������B�����>��qn��c�!r��]WU,�7��t3^�[}Egtޜôa\����M��0
X ���k1ՓG���Ne���jV888�KS�;k<IQ��p��*
�Y����d �!��������X�>����J-}M��ЉnaJ;�*p�}�HS���%:ւۍ�h����&��ft4x�}�Af�Q����)y�Y'����l|�T��С�B��i���]J�8k��HVW!��,	�50��Fg@c�� 반���Ub]m��@��Z:��I
��E_���sF����1��P�#�B4R.G�
Q���ȭ�a�M3�	��P�XS-��9Z��d�-oSX��	���3#��5Q]t��fUP�I�i0p�5�G!Us
�v����H��ʉbB<��{�B�끢|R�W���K�9P,�5!��^���������q ���ȓ���`�@L&����xjZ��8ͬHW�� D�����W�6կ%�P�a¥��6�� ;�iMh�;=}����A���R ;�2T#������9�X�����`��)�RۯU;����!�QMFP��U�֜@z�2T��|�z�b[��a?��Vy�JP%̰z�\,�}�̡~�@���hnH������xAAjulC�c�g�a��Ű-q�1�j��M�{S)�>��7�Wy��%�&�h����C��0N4���;e�OT�1�[q�;wU�S���v�N�s_�P>ȥ]��Ꭰ�˦�4m�R���4#1�Uz�}�u� D[ys�v�G���!.(����'	�74�_$)�����������}��*�X�|.�'쫇7^��l��(rW%�'�L}C��I�u��LmJ�4bd����u�(��tx*\�_]o$eׅդ@^� �Dw=F#|]qyy���NѨ�o8gxv���*z֐}SR�ʀCWR��F�]֢��Ϛz�3, '�-����\
��BS�x ��gr�����4R�P��zʏQ�x��fG����ɂ#r K��0��w[t#����t�ȝ%$�nr)ߙ~Qֳ�HP�7�����p�D�1�F���s�S*X��E�P�#E\��?�$�*�4
��M���{w_RF�ldM���\D�v�y�^#�V҆ `�d��_�O��

��V�.�XJg8}�q��vAAc�Q1<>:��p�ֱ��h�8�5����z����M?y�w�sПm��;����3,�c���$%F� %_�!Aǈ��dJ4���ᩣ�7�2�x�g0:�U:�
l��Q�@���a��kU�&���Mq>6���l����Y���<A�ű�VU	G�E�2f� ���}�{%q�.j��2����9�eh$��R���v;ܨش�'����:%Vj�4>�a���L`Q+53"�B��~s��b���S��t�
1�a#N�?�/\
�!L)k���9��A�Ջ���쯶��f�Q�S��XJ�b(�3�tD�[�
Bd����:�n����!�X�"��h	B�ku[��7�:���<����셧wX3(=�ERgr��c�@9�c�T�dU_M�\[�Ƭ���uҟ���e���c-��q����azy�8�$���WϾX71p,\yV��T(7��Dz᫋/��ց����n�;��;?���~W�<�����N*=��_�EŚ�7��U�I�@�UT�LS�uFn��{�����6�}Kz=8妦��U�(��Eƚd��"�@>bq��q�(�-�)'��<_�>9���"�Q�㏒�	l�C|�5��ejh��t
$�t����rX�[9�E�����uBs��OgtQl�n
��L������~�T&%�ה *�H��;e*�XM�c��hJӷ���u�����27�����Z8�x��%E��~3ҐH�Y��(��f�D5\j�G;f7��+8�qe	o�_���!9���?��ZHƮ�t����tt�ŽX�*"��y2�]������SWz5����t��g�(�����k\R�K�Ω��-�ӡ(�������U����P|S�����-����WF�D�g~?��wc�����B�ӳ��y<ܓ��N;�Vi`D�������C��^�`�Z��Qt����1/=H��jn���x�ҁp>���1�,�w%Y�u��?ǔd.��a~+ZY����30��	�?����N�!�͎vkGP�HH�
��̭��m��p��&�p�Ӯ/p�q��ia�UPv���!�r�mU� �(�0n�Я\�m�w�+�����-�;_��VGr�ݘ�u+.M�P����S2�
����CկW���
�Ʋn!�$0�şH\)��X�j&v[<�_�W{�p2���2g���p��f�~T����1+�)ſ��ǋ��e�'�,OBr�dZ�M�����+z�<��^���54�1;b:��Zm���])��>��}��V�x�uaLğw�x�D5f������l=˃�lS�1��wKie�ɫ�zH1Y���^C��B�IG{���S�8{�g�-Л�"������1�&�NMxZ���>
�m5IC���Mo�ٮ+yw4u�.zSF[���a�R�6�N��I�Y{_���O[�=�^�z��Gqct�Y�1U@ι��MG*oGIb��V��� J�L}m�gmx�XL0	��ܼ�J�Ƴd��U˽��S�6��ql>~������c�Z�Z��0/Фne�Rlz���.X�Ś2�ڧ�34Q�G�t1�dZ����ܰꔈԛ��l�W���g��e�k#�~�Qi�N0͕h�10��.�a�oE���C<��L<og��U��
�Y�2���"z�a������=)ڜX��gi�Da�a��iN��!O\Ѭ���������[|�`�I(J���a䂐�����
(�T�,2���<�$����rAI.�W��`q*Փ�Q��f1��1CX��W��F$- z��R;D������m�ɼ�����%�_FGO�w�l~�G8��I�	�}����k/y��m�+�PT-�|��ͼ�<p�0�o�hI7ujB���h3'C��r�P�R��U0
"ZY�u���Un�Ր�ݫ��p���͌bpa>$=&7�5C���Yn%�Ң(�XiV1'5��	��`z"bc��������@X�<�.r�+?�[עCh@g�����Y ��gFY(�/yX�����DXՊ]2��;�r��tG������������Y�:->{� ۡ��'07[�k��d�N%./�0L���0PʬmS�!:Yl&�����V��h7�����$�CO��y�.[�h����|�ӿ���S�sҖ��"��'��U0������YT1㒴.8�� ��vi��pLA5�[ueC��'C�fV�Bl}�Q>vwA���-Ϲ��0��`�*��x�Ml�6 ןD��D��i�ϙ�=� ����2O��7b��1t�����<.;�3T�+l��>1�*$�>�Ⱦ��kǗv9�)�Gn��h;��t����c�sڡ%6mE���ۆR\�9%�4��]���;�I�nc���aRh�wo2��UG|<��#�rQKXC��)Ɓ�K��Vu�rl��Z;J�b:U���&.ݳBJ]�/�U]��	����������m�7�E����^�Yw�3<?�޴⣫�[�yꝌ2{�/��J�uPx��s�V��sas�䷜A�,ć�:2lD%s����g�]�m�m�D��e|s�_ӯ���'��6O��{K@��=U���5�	jw	�;�NϯR��Z�>C�����Z��o�F�]�L�c/�d��ܫ�%��)�A?t�N>;�"e<� 7g��T������}H��Z�X������E��y^���;�b���,}
�kA�$Uh�}/�_1F����kj�Ǔ�� Cx�g�\E,p(Mn���Gi�)��>��(�步���y��*˵�9�S
�����������B�����o�0�Ez&�R0𡇃�xWZ� ����m��gw_���<(;������k�CI����(��G��	�,��"M���t���"�.	b��:>�c��\�}!�7HbVzƋj(�}�J��\>ACI��߄���Fm�V���q��߂�1#��z�����?HT�t$ �?��"W6���������B���U
��[ �e`ɣ���zn�٥/BPzgyu�?3r &�}��*`�d���W�!ܞ4m�����$�'*O�
��Q�s�I��T�9�f��1������ـ03��ƛ{�|1&<��{��-�nW3�;����[zYE�m�����	X�!��,&z�'t�X4��{.����Pr��Y���럐G��5n�u����&���2G'�lbAt��-����x�>���꿾��ZeU��ٺ�C�_+�֚�w��`���\�q(�2LL<�t�*1��-*>s�ߩ��7�ը[�q���Q{bL��}+ݥ����a��TI!��)g�;L�w�{Ƽ�qʃ2�|�˛a�ClN7�����5�3ݟ����R�ۄ1a��w�7XD����6JQ49�~	q�J���-�w�I	U̔���Q�GF�5��{���AJuF��A-B��E1��-.��EQ"����/����U������N�,_j���K�Q&A��%_��oۼj`L �|zDO���t�h�n_ڳ�Z��FsB�~��Z�7�R�Eh-r!g�eV0?m�Q^Ej����}���k�x�EgT庀V�`��^�"F�h��QB������t1?]=?I)%��E����5\_�;�Ă�Ri��ǦN�f2�[c�U1gAz��4�m�7P|��������g&���M�f
ާyP��M�k�0��8�a%��bP����A#��e"��ȡ4	�� g�m���̱�}��L���n�L��u7�/J:� 6���Ѐ���?�-$Aq�Kd��q�O�s���H���i����F�F����j�)i�������ea�&��˩b�Nhj�?+T�
~zL<�;���� \=Gf�\�c�V}��������R�n.(�D΄�C�
��#`<�RA\��<*41��'�W���A��c���w�$�e�9�\���9A\�T:�O�,�L��/���(J&\�}~���;� ۜ��n�A�I�Fe�A8,�4-�E��Q�� s����o��qJ3^��wvOw>"
p@�G�/lnW��S\S��(�����qW��1������3���zH��쑁�[�u�R�I�1�{f�)bd�]�LIO +�[���*��)a]\�I��vdľ�q̛��縓�:񏕟�1�+�)uRY��~sh�� ��H��}��p�$�l����2�����(DB{^Z��AL�[�3��7JŻG"S?���%�TSum�i�jp�$�f��
�U\p�
X��LA?ITTh\K(���:�iY[�MG�ǻR̬}k��&�zU��
��uAs <R�&��<sR�����������:XS�|�u���e��3_ !�g���j�h[�6椢��%F����<��@��W
`>X��[B�4b���y<o��?b�V�<&m{*'���#�����)g���;?,��1X���*4��;7k�[}ᰰ��&[�g	���Ճ��b�H�zmI6�.:�v��;�3@��s.� nI7�?����HEp#.���ͩ��V�c{�lM��*�ķ�Kk�F�3�(���^�
���^�ԬNџ���-�������4�vk�LIdaUqϝ3�8ټM~�[WI�b���d������[�Q���3z�U�m럨M�����b&��Q���l�_�ә��ꩥ&^���K�N
K�V_�2R�H��^F�iP�@�&څo\�*'_��6F�W���ZQ�;Z�L������J��b8��[c ��g ��:u����=�*-"J�oG���[�.D�$���~��5Qd2^j���� `����'�I�KQѴ4x����>��05,$���K&����A��kBhL�M���������A�'����K?���HP>R�KFҊ��X��4��,�3��zZ��SF%�G�Xro٘�����#nM��ՙ����)�Ζ/�`�=9O�N����� ��έ����5��
�B,'�j��4�4n�_�o�W�- �a�����i�7;���ϧ";��&��7�Qڒ�F/kTj��6E�N�R���y���7�}0e���i�i?G-��C��^|��ev��}����Z}�	�ݹ@i�%nw�,�#2��� ��k��L��l(����P(����K�ܳ�X	z"r�2���D��m��-p�������Z0�4�6�U�8�R��w-�}�@i�m7�$�d��UOW��xM�{��.���?j�f��G͈|�f�q��n6��	�A��v5 �J���
Gf	j-_��v������IV��"Q�>��%��QçAҒ	�m$7_:������`3��ƭ?Z)5L�Ā�)qH��ދ�hS�8�X�y����JAݡI4,)��L�9�q�j�,�1��r#U����Uv��*\�{\�:�p#G#C�QB�Tk�6�y �+Ic�s�QDU͆�bi��g:�Bk_4�BΣ����&7���$+�P�wG�N�ì ��@��3�$c�7�:q��ˣMW;,�E �g4z��cϊ�T�eG�Q��j$<�e�kzX�DP���5	�o�׶�Z�����j�����y8R��s��w6Esb-�@5��&\kȠ�S�r< ��j���,����'S8y����8�Ҫ"ݳ���1�
讏Ն�5J����~��`[��w���{1�=s�������;7�"<Y;��V-zZ��!b�%,س��S�n:�,��̸�G�`fǮa`s�¡6���)�PPI��q$�b�����F<�����Jv쵅��Je$>�ӓ\�7wWǨ�E"=���퇟^x�5Z|�l�XM�@耙4���wRD��f1�����Dֵ�cr��G��8�<�j���͔�������.�k[���+M�i�(E_�(i�fc�7|q��i��*�mYkY@����}`�b�!6n�0�/�Ŧ=��@�f�����z �<�_Ye>�<�QRФ�q[9��M�1��N���o��0��&J ���j�
T��Q�1��<��.�hG��'$�� ��\�q�{��Q�N����MP�K�C�o���~�bջL乱�wȧH�C����`�m�Ms�G5������`���Ȗ�й`Ȭ���[[���8��>:��*��c*e�� �wBs<�J�j�`;�d]��y��c��fx�Qʜd�	�S1m����Qs<��:�w�p���o]zr�&��aU<�DZ&y�l����c�!h|���"��C5�
��4\ߕ8,��h���	��=���`���+I�z;2����:���z���:��N_�i�M2�eR���&��=��ų�j�)��ɚ:�ۃ�]����Xd� �D�����E榥^��*Mt3MR�،�I��!�TSW�@'�f��M��	��ޛ�+���-p���#�2iy�'(>��Q����eJhu��	�o�WC�A�gi��H�ָ�/F�u�?�����-�+	N;�d䛑yK֎7�M[F8�#S:A� ԻP��h��̙��?��*��+1�u�#���c���kX����hL���~��)��ap�v���4H,�L�H� ?��s6� E�@-@Ib���ܰ���WV�c�Z�-.��b@)��T(�>6
x#O��Pv�a������ݐf�Д���J�},>�q��nb�\�#��Z���#�J+���Nną��a\W_�	��U��	<���'O-���>a�q��Q�;)���]X7�I� �b;u�V� ���K�Ru�pâG�(�(�u�2 ��˞k���0'���={�n��xbď���9�nKZ-p���Z,��f>7uX�qxB9�f����яyb$��b�������Y!�C| ���
|��J4g$r�:�o���3�s�<;�Aw3��P�)D\�ӟ�w�n�=4���w�*h��R����+��_�_iH��ZJ��d˲������M��a�r�J�+�eEȆ�֘���-V�L�%�Zi�X���x��=H�	(���7�H�'/7l�������={l�_@�V��'��6d�F桺ב���+A����518�x[*$���|�
q�!Z����}�I�0��
�Z؉w�B�+jk2��,OC.�~_������Eo
�'��A�A�7�C�HK��Tػ̅�>7^��HB��y;���9� ��	���1G��j�3�N�?଻xF.��,��L��/C� L��CIȏW)��󧾾BςA�r {$SZ.�>m�oh�og��)p��VDNњ���;/�B�����9)J�3µd_��R�y#U$7TǑui��V���z�ҰR/���m��G��A ����ك��d��b�4�O���ο5	�8�֩߳�p��@�A�q3��y���f�$P�����H�VϑZc����3-�z8�+!יf���D�����f���w��fy�S����n��i�e��Ŏb�1�X�)���u2�*O��Ϝ(��x�N�`���s��M�0wP�պ��m��L�[�,"�k�W��x}��$_��H�w�B����w��(?*�7]��%ݿ�-��H,dU���j��D�������V:MBĵdV$��z�8v�kh-ހ}Tٗ�(>+<�4.���B#���l/l����X�~"��p��(��n�;\�ě�q���T�Zt"C(0g�j��U��ę�7�'�_��
�|�"���,B��ē!B��<�Vr�+nf.N*�6v~G�{!	2�����r�����|;�i�-�4#�zB���dw��v-2�{�T��g�l�I$C;��$���6ν.�4ޠQ��c"��2�!b��:Jt�=±�)�t�	ѮQ����6ɛ���0Wp�i���� ���fMM�o'W�aŬ�{pD_y�x�?���:.p�͋�G�&0o�z?�0�_Ҝ&����R||c1B]��W�
!?���LO%�G�H ��ד��x�_�A�nȔ�@��p^���`P\E��}l08^=��*�������3�n�]��h�T$�9^��E���)��A�<M{�I�*�S�b�7�,6���b�!2#>��`��<RS�
%��Yy�<e�8�YEq�,� ��@u(��䍍3# :aR�[à�ɻ��1865~���³�sO���g9��i)P��"�t��چ��	��Z��0��+)8Xe��C.�'�"Y;Y@?s3u�H4$�'}�� �R�[!m�r�L�L�22Ơ%G�^K�3�`���B�\��M?���gӰ$l.�;��Iv�|��Tc�C�V. �2 صt7��Q?��)�x�n�z��`s{p�9�؜��o�E�F�Y��6�'n�^h&��I�e8A�R���M�@L��!2�"����������{&��Yo<�9��A�����0�T�Qh���{S�7�:��vY{��������������As�d��o�<�֚�Lۉ���@T#B\^|���uԬ��#/5�;x�Q�_�/9��,#K�&�	�#�[�Z׷�kͤ[���/���Z(��EwU� ��_V������<�S�E����hh���r�L�*:���
����OR�)�4Q����6�¥��%�K`�4�ab���3�fL����Jc�t�J3�>xI+�]��SAJ��c%�F�uv���>���I���c:ع�*) ���Ӌ!c���N�h�"G����kbzt*�\��"�$��9L�i��sq>(��D;���4��ē3�Y�#4<��!�tl�I��¾����4��+��~�[K�d�;�	0[��Fb�Ѣ��)c)SQ̹�etZ���q8�%&`{��C���R.J�yd2�'1;p�������؜�K*�P0�Tw��-����Q�h�Xe(w
�{���
�:,q�������>�0W>̰��r�JB
�З��pI�6.�ъ�W�}J�>�n<Ųyn^����r����Fl%�Z�9�ec����(��]U1�6����wưI�/�2kKe�t��VE��V� /�0����&�'�j��Tn�N��,ʿT�9Ꝓc�HNn�@7@?:�8�<������u�-�s�P�+�Ӎ���<Vɢ1'���}PU8�G@}dX��C,49��t��Z��)�(>y�6=*�4b:�{'?a��@?�[�J�wl���{;5J\<��(`r��!�E�LgP~����!bt�8d��*�� ��*u�M�/>���wu��,�d [2�u˭�����^���5���B�Ӹ����9�S�#�{cJ��
]�f�k�܂�$�`�% xr����B�`��s��Y�R����ڜlT�]�\�M58��EG���P�V��N��~IS���Y���I��TV�*%i�I]�;l��p���O�KV��v�Mڥ�ޭDT��	�0m#��'T��(��`�1��V�y��
�����׷gk���.�xA�h��L�G(Gof�0��O_�C	��L�%��@(��"S��mB�Ej$�Ȝp[n�7V��9I��钇�Ĭ�"S��Ċ�?$�onPI]�^�ьW)OBjNi~JU��H�Zh����Ob+��l�np�G׆ !����_b7G !��.�o�[��fFP��8�&ڙJ~�&��z��?ֺ
���1O����$� ��'iJ������;|}ux��߇?�"�z��S��@:��h�pI�äZr"ɛp��L�Xc�O �wI%��& �=rR�@SG+��[+�7-c�Q��Z� u%Ou�S{ٌ��;q���  �d%P���av�XHp-�b�nf5�3Q�����u���ϐ�V:|��JP��b΋\ Kk�<j�Bl)���U����
05���9Y��A�<`�Y��9?]zA� �5�h��2��0�I�?��Y�3���y�Y2�]��^'�.K�K�*j���*��֜��$����C+�C\0�V�*�a{v���F��1���lk?]�L���	~ v��}"H�m9������.-�����<�";��ÁA g������&C >����g��9�w���N�D�߰z�0�pP�8Q	��vs���Ci�(!�2�	Tp�9�d�F0+n�W�J�H�p�ʟdo�����eն
�{D_*s�FoW(E��9�p{X��#�&Ob$��	����;8�fc�6>�$^�����J5ϵ=hT�|����)39��ZX�Y��^��ʻF׼��^��Ĩi9gM�M :��S�h�+Ɉ����p��>���яBX,4\&�a�e�,�:�|�p	ЗjZ?	6��X�#�Jg]d���߲��K�]��Ml��=	P�B������ٝ�,t1G�Vqf���*�I��!��S����,.�_�/��m��nsʙ_�;�k��[���O�Q��A���r6o�KD��z[�2�}��j��3dY�*q]�]/�~ ���1���7��YD��+wY>5I>$��UP����uDdP��\��2����D�r
�߼�DZ��?4DY��s{]�ʙ��ϊܷ��e���3��8`-��vS�w�(��^|��?��_��aR���o���?��W{pI����CvK�QM����o!�愦u&�v���[�Zf$,���Os9��-n�����������J��<{5�!.����o�p|W���)�4���?lX[�~&�Y_��4a�@+���g��/��e�X��0��y�Q��J3	ߓy8>��x��zC}�X��^
�H�����
U�T[��ØP�NE��N��mF��{5@VȐ�Ҝ6
�߄��41k"�/�;H��+�����I�D��TO��6^�)����=�e�+����~�l��k�ǩS���#w N��zhl���O�~��T����ԆT�`Y��-�H�6����Ӊ�vsҊ��67�?r�&�]�qZ�a�3%|���`󝥴�0�qT�d�Q��-�����ؠw�=W�(
�]F�'?�;�f��C�2����ƶ�P���'bA��ʦ-zrRe�\^h<d{x��P�����4fr8�ٙ�&�#֞��i�^e1��;w��9q�]�@ꊲ�)��r��.�i�!�h;.��Ɍ�*�R'���&����v��Ʒ����G�\T�W_�䞔�G���]C��Y���x���/�J����Q�Y���b�l�g�t<��f��	��7�]WC\��giȋ"�͐C��7��!����ܸ��t*j&��T��p�	��zV6��#����e�����f����$�Tg
*�؏����tp��T~wᩤ��mM�w��.zȋ"$��蘹�}(]
.�j��?w9%�����Z�a����҂/J�66�o��9u��9`���{����k�X�خSp�\}���˳�v���>�$d�F�t�*������G�=ȟ-�/ �!�xG�+��g���Rbb!U�����@�ݓz�A1N)"����ms'-䶈,�����C��i��B��y��0��}�AGC?yT��.K����k����u�m�4�	��~���^�qv�ʯ,�`'$Y� ˈn"�Y��}BjQ,�'(�f�+���@�֏m^����J߈�l�2Վ��0��[ �D"���5&+|2���+ղ�Ӎ)���u��,"zu���k�&�I�KV%�(WBbz����ΏJy�L95A�?4{T��*�'l���i\o��	��#C[k��N�$J)Z���F&MͬX��q���>:�/��j^_����U��o�@eץac���)C��v$$1�I��N=�g-u�L���+���,Nx�p�ej���'aI������r_>�E�Eެ�թO�K=�}����v,�w���&-���(�>Q�Y;h�y�n�B,�E��;�U�xI�\�q�����&�S������&&JgT�x�kc@����Fl'���k{ 1��#Ej�4�ς;W� ��C������:���A�}1n�Ħa��߆_�n<���E�L�x_��$,f��
y`�M��(�ۯ�ŌV��u1�.���C�Z�ی�xpW�ԛG��*��aGz�ʉ���R�]x�"�-���f"��r������3H3'ʩ��dW/���DQ"�y,	����=Ě�7~��ٍ_�^���^�\�fa��2.@����B�>�^���5�G�b,n�d��r�c6x;
	�|D&L �R�,
��N��v�����3(��B��+l���M?̽ےP����A}&�Nʅ��7��ΏB�Tp_1�S�wӚš���M�NJ�)QFL�7�4�����Zn=& �%�]��tX5'%/�c�Pl����3M��P��@���dKn�Z���g9*d��?�S>�����X��l�7����c~c�S�-����+�m��t�4����?S�z���.ߢ%�~2B�i̿w����?X��5(^���`�&���)�n^e�4���H����6!��
if�˞-�7�q^���, ����a���;�+E��qj��D%��a��ăN��rG�T�B�hK���j�E�/�Ȭ,��r��>d�����`��~^�����-�U���k��x��`����
|�C�����4N\X��'h;�0%����`\.e�ɹ��q�ޫv�S��9�V�x�-�0�y� d	g������dk6md7)��s�4%�$>���|�dp,�Q1�*ZUU��P*��򭳍TT��na�?gI#�VCdwE��,��hZ�Z��W�5�KJ����I��>���Uadǿ��q���_��E���6�FL����b9��A���&=�Z�C���b9�J74ԍ��IsUR��Ӄ���\�D��]
�!��b������ ��dق����e̙�'���@���u��ɷF�>���"��4GpP�����,��rÐ0�S��Ya~l�8���!9��f�fIB��9X�źH[�	{�[�T�ȑ:�����P`��0Kn�r��) h�M��f�4g�@�)L�VT�\:-�na�4��8�Ϝ���o%�m�����:-��=�9w���po } �@�M�4Re�}Y�����5�P���KA�����*�1�\�Ԯ�HR]^�-؎���.�F�����a�C�U�,����"xU�QlM�Tf��i4⣏��˘'!����ܱa��w��}^b�i��у��K�KӅ?�{�bۉ��q$�s�>Ph`���i1���R���{��Q"��y�����	T�%z8�ݿ��0m��	j��lě��&��Ͼ"�#	E�yRz�_P�r�)����� �����U����)�[�\X3��^V�8��ׄQ�m��%{+�!�/��(���,�8�V�L����yɖ��H&�{��t�q����OO�YyR�~�1�ID�������%Y����!3���r��hΪp˅jA6R���g���"$=��1�u:P��<�ν�xWV�O�p/������J��Q���c�2w:P`P#Y� �)�f�# ��d.����D��n�;�G�9�n�2f�KD��|*�MmwҠ�c�2���P3����h�7��� ��s5�;"Y��l	�^����b��#>��B�Sj0��Fi6�����*۳da��ȗB����i�8WܯJ�rQS 4h+�lס�,y�Ă7DcQ�|�$V��o\V޷G����ƪ�p���&��s#�!r�]��r��nh���51�V�[�
 ۜ��"B�]�K(t8r�X�t���'��9D� �	`~�l��ul\H��~��5��k\�3)$�I����� ��}�Z�z�t��������j��n?��#����G�
Oۊ�P���:�v-b�B\���K9�3_�9˪+�xV�#�T������.�������Js�y��Ke�5�1�P�3�92�3�U���/b�%��N�0%�_�A}��@ֳN;�7��Y��"�>�.�Y�؅^���GSy�|8�!=��cɁxi���)dVcq���������B@�E&T�>(���m+=x�Ŋ�v/G�7#���%����8@!��.�ʗ�Σ�V6CѺ�Y�w���u���r7̏-Gt�zY�:&3ͨ�II۪#>(k
"���e�*!"�ג�x�7��@But���d���jH*�}{�����>��C�?E�%��e��癏&D�S~�}t���n�$E�+��W�J�� �(/�YҡtSL|j9yCk�/*�/�o�؎�#I�l�l����F�-�~%=��)�$Ǽ�o9\p�5�G�v��vSh
������)
��tEgg��fbj�w���%T���������ș{���ET��rG�`7�Ҕ2�=>��X_n&�ֳR�����tv��>֘ģG�!k�� �?����)"X�4ȸKR���x�D쯥M	�,ܩ�r�+CuD�!^gԉ�NIj������P�����Ҿ�U����Tg5*;�,�C�!�i�%��\��EXG�I-�s���Ł��@оZ��kW*qhَ�A��)�o	�.~�bu�\��vF>'�"��RQ&����<��#��8(������YV�F�@��T!�)�S�I53�G6&��e�j���,{1�I�N8���)#r\VǕ�U�$�-}:��5J��d���pM�A���kp������M{^��y.&p�ǒ������\��<�ut��B_Zw���y�b����8eW%:=�oY�7�zQn��yσk���4�I�v��zbI�<e*�]�
SG`��%<F-S��1+����XW!�eo��{��>�9��}K�V=:31�{�nd������o�%�>:4��A"��R�'�\��Ȳhv�)�5����G�X�g����_#�`Y��S(�eL[��r�3c���=۪qU	0q�+�F�G�y莵-9|5�F���;a#�A��O��������􏎱��[���JH!iDn1&�����kthY��A|�t��Cm��U���m�!r�^P#Q�Q�u��B����f�iH<�� 
��ɫx�hv��g�L��(�TV�t#q���C�8r����J$~� ��[��m�P���}�g�d`q	*�@�:z݋���Dʲ�Lb�	��J�u�E�Y��m���E�F�Y��V���q�n����S��ƛ���D�i��яn����ɮ,�b�.��1T���⌕ְ1U{�?˃\���Wq��~f#�%k��n
zmB���n�ڛ�j�9�=�R���d�dF��k���~��K�Xd����������x}lj��tU7̏|�w�~ŬwO:�~�<�98joa�^�8�:����@Q�V��O���=I�B���/���a?>g�SQ��/�f���[8���� *Ldw��x��G�*�����,�����K ��5�֦J��$~Ҷ�&֝XH�d�v�&y��ߌ��`@Nӻ��^�U�Zx�ؠM��D���ĢywP��2�ߡ}�1aPV����R�R��F<xD34�������ӕ���4k^�⑴�1���v��F"NnWMizo�n��x�P�
��]o����x\vw[�n�,�](@��~"���\���[�H9Yî�JXJ��}|�/of,M֙�M���L�W���@��A,�Az|T�U�\')mR ��ޣ4�!q����4�bsէ�ol%c�2+�O��X�j�+�2B��2x��'�l�e��{6�s|�p�I��Q�S$�5)"�\n��Ĳf���'��nJ!�;�� aG:��RD=����@CmT��q���2i .&����\��";c�����׬M;[]�KM=�i�[�{��W��٤��N��Ӂ���A!�6�6�� C,�x���d�`�H9��Q�-=٫Gb�4�r�'!�4���M@�T>��V�j�G-�BY׺�|i�b��}&� {بP.Q��}�I'7q ��CvX3�W�O��~q�˔B��64]z	2��؀�١�8Q�D�1�4�L`w�P�0\�7�6�R�h�څ��R6� ]
UpħH�pN���Ά�m�4��В������@~~��i5�P�aYy�	��SӍ10�[��{�t-���9�稁;���f���0�$�Pv���֓Tʪo|����]S!G�W��M>s^f�OH�x��6%�����'�Y���x��R!��Ŀ$���3bD�Q0G+��@11���-�Ɏ���Fp~M5�I]\�#ib����}�����Ʉoc�6w/�yv����P�b�M�wL�<���{S�8���H��P\0]@�ݨ¦\� '�&w�&�09�ӱ7�s��he�fZj�[m,W��;��rߠy|���I�&15���4J���'4�D�L>���A5�F���Zo�v�'�pd�\���U��rj.�U�M�R!�8�u]T�?d�ad�<����3KH�	���G���J9P6%ڝ�j}�+x* ��MO+�di� њ�Ť�I���O5��̓1����W�����;�,e˝��g�"��l�lh��ɵ��ɜ����Sy1�����$�޸*�i����Y�/b"���$YW�!=\�cV��^@�}8�k�6�<������[ޠ��V�ɖJe��'�d�ڊzB�����(���+���WsК�kC�H�r�{+PX�jx���j���t;���[��q���ɿ�t�`e��o�c�����]���|���׼����,�č]~O�R&>�.�ɛ<�$� E:%#B �Eׂ��Xy���F%�Ų�����P;�M�~��L���𡳛k�-�o��]T8��JE�x��D��O(�K��Z6�6�J�w�"~���˝���(��Hx���{_��ìy���)1�H�ؗ�bI=%�U�h�D��*��%�0�ӻr�2e�c[�+��-�ie�K���7M�QBI�D^�{���9��L'�=�3�9��E�J�S��[qJ|��gKH��'ҟ��TÇ��l�v�R�4�JHã�-]�k���b���G���9(5���K�6��1�Е��R7o��"���9$\]�$1����t��)��F���c�RR��|p6Ϧ�Z˝� [-�=cn<_�&����y$�Z���)-c�v�l$�RO;�c�t�3d��LN>�.Uk���u��<�	��nH�s�AR:e���+1D?E�N���Sv�E�P��(}��x���b�v�H$�p	[�7�>8�h����$Z�U�6�8��8��s�5wS�i熔U��v��K�_P,GG�Ѱ��D>�S���jm������E����,�xORa�&i(^�yr��9Ὼ.�����YNro��uZ���:Qg���e��:-��!��0U�N�ϵ���dWWn��z�v֎����\�)�ٲ|G
�����a��?�j��ڋ MrW�����c�z��GӲ�o)�"�u"����N50_�>m�	�jѭ�KY�P��"_��;K	���u�q��t�_���7�
���9�\.j�`{���h�7��<C�l��0y�����W4��aZ��F>��F�4ƺ�f���L\���W`��lNPd'��#�4��%j"]���`Ͼ-�{�i2�Zܽ���<K���y8��i�`�JZE
Y�!�/�#l�A��gF��Ꚛ��jxҏ�0!d�V�X�1=��}��Ұ/�o�$��b&C�����p����X@�:�e�(&�o�+�Nu�l��^j-Q,&w����Z�].��9�1���l�z�����CԿ����5y�c��[�f�U�+ـ	���E�����>�¼��kݖro0đ���փR�I>��:��J!�����Z�Α��O%)�&�M��:�Ұ��W�������S���J��������zy�Vqi��"���R�V�ԋ�¼]��ԧS"��-�hW�]z�&գe�j B_#�����B� �Y\@Gۏ·F�h�{���6��w~����b1lߜRn�ъ��*�I��Įv�kq��س+�J��|�v7������+�3e7� ������q�E��T�Lp�
���5�z�F��H �<�vJ�52��`���NF��J��Ԯ}��K^��*\ci��u�7E��ϡ%�bh�#���D���^��zh���ž�̢j�iK�d�\�I{�rLp&����"�@ �x��2bA{ ?(��]nÀ�f��EE �d���]��W5��da$��;0<V&����^�֝���Wy�Q7�����K1��iu	~e��XL&��TH\��F�*s�q��q)P��f�&���ϕ<3���<i���>��$^s��P�"�T_�9����Y����%G1'M9�!�)���S��t��m��k��#����&��,|RS3�&�g��:D\�}`��"�ˈi�^_��B�*��M~a~�p�  �����7��V.f3!D��'�#�d���M #��AV3��ƾ�S�A_a������l:1N[�RZAd�0�b������
[@���j�0��yw��[��}��mn�T��$0C�L�'ϴ��{�o����(͔��o����!�T7��'�U,c�î��1���.�0IT+--�'���FX�{y7^7]�qbR�h"Ϟ�7î|���o��Ξ5�(��p���3�]	v��0�ԯ�3� �z�caÃ+��팰�m��i�f���Q1���H@�'{�bZ��7P%ߝ#�6�D<����I�F��*�0O�;>ٌV��T�N�&���
Y��N����X�]MEn�۽M�!�i�;�OJ�t���O��<�|T_N��p�z�쓘�*��</�$.A�'o ��Z�"�W�ۢ�=�X���>r4� H��Wt&�#B�	W�y��W�բ�`��Y�/3~���-@�N�5.�E�R�����j꼷��0�$�;Z��G󵍙�A����xQ5�g:ԋ�����)���t��|�W��_!*iH���L�8�+��)��2�y~�3���rѤ�I���4�N�\��d�N���}���[�#qҦ2Nؕ�� ��#�/�E�ToՐ�V趄%t}��Y(DQ��00i��M�R��s�l	Y!MM	�'��w�?��Z'�V�,w�SH��I�ܑ�G-�;��������1��	�,�iDTG�3�pJ[��r{��0
�`9�V�"����p-��Q.�wU�7�n���[$@��?1�1%U>�� �����J����,N�f��_� + x蚋L��3T�=:�GZK�7HF7�MlAu��Ÿ�����0��@C"A������ Sz���"'��Y��D�����s�@՚ �뛫S§�o�Ee��v&�1 >��x�־��k�2zyF�M"_@�"F��s3��d�-=��̮3�]	p�Ӳ]�8��`�����F���X2-�R�;�ʃi���H��q&~Χj�@�s3�:�B�C3V���:�\����!�7Q�u�4����2j ?�~!<�I�'��۽f{�s5�q�� �Ω����z7q�3���yw�]5?�\,�']S��v�{[v9��!�U;��Ղ�He����<>�E{�/e�K��	���BJ(H���;O��,[AWn��5��Ek詝�J���$�=�/)����6f���9���_Mj�+埐�Ѓ� �i*����AV,\Vz2�S��v����hI�� Uq�<3�Ǫ�wx����QD����e���ڙ?��jE��CnZO:�b�ܤ����<(.�+��d���ߟy�y�z-�*�.:b-	d&�bG{_0�a��2�7H�>zlA���b�sh�W
�"�47ωq/N$�Z�,\�ĕǛA�����-9��όX� 1N(��j��3���,�1�&D+���G�)��Bz��_�h�/�@\d%���@������8ɑ��Zu�c�V�6��r<�5��Ll���L�����/����XP�[���>".�<
3:�k��˫��^k"����k^2�v+Pt�.;D���;�-��m�g=����D�3E-d��NC
Ϋ&F����Ul�I;���S�����Om
��Ȃ�s�k:fS���>�F�+yd��w\[@��x�5���m#�^n 	xd,"։X^����i{u2t�E>�vm�&ZmB��+T��=`5:����Kԕ�&�5�~	Y�R=d�2���=�S��0������5	�Zav`ɪ�J,i����d�������v����m.��$������Uow�%wq�E�p�8m#g�iV4{���TØ�U�l\o
�?�	�Fsά͢����S�hQ5 �����,�:�;�m��Q���LI3�Tknտ�ā����W�m y�*2T�q`\�wgi�د.�eZ<�*�x�>�qgN;E�<	�����vx����%̉3U�t�Tgc�|!h����Q=��CCب�����ع^b�X���0��{��6�c9!�mҡ��D�Q�G�mC�P���32�8���!%Hns�HoK;x�Z`�M ��f�ct�a;�!_�M��{�gꇅ�FI~��F��k��&�>k"��������	 ��w��h�3b�1SN��0w{&���}eUf������xO�%��+Y��� �M�����V���3�����1�G*P�?����Y^kG�J������>�-���	���'����{L�{*aխDgS.��V�ȹt�v�VG�>�x暑�h�� �G�2b<b]������ �{����U����9��g����hɵg3���%0�y�ƹ׫�+_{?����Q���m��?���1dy����Y�j���������r�é��1��O�X!/* �Z�����ן�Xis%Ռ�
B62�|֟��q�=O�G�+���ƫ3�4�n��k���8������y���ֵ܄Ȗ��دr�YQ����T�7˧0q�,�Ӄ�&��O��7Hqݰ剜x{M}*�`��+
|��f+�ކs��R>��]�"��CV���?{d=S��HT���6̞A'�-*��@�B�R��
�jUvh��'�W��Ə�ę��ƻ�e'��6��/PJ�r���G?K�l��+��!)��
�S���)oPo4ɳX�Un�qS���AG\�B�Z�Ƕ���afV��OI0��)�c���Քt6��\�Y����3�ָl�B_?��r>���S�2�C4=  �a�q�Wo�D
/���?;��b� \|��a�Z��
9�"���D&BR�.���T�R���נA`.�a��Ĭ��
�ݴ���Y{��eޖ�Æ^!���iF��$�e�E<�"����g�q/�n�!* 0c66If�\ ��=ʈ�A�Qp���M�,��C,&�P&8抗D�,��g�A
:�j�t��~>���
B�2sF��&���{` �N>+泪�����t�_E`�܂������WB�!dNp�6��"��ҺE�bP�F=��.'��Xg���d#�7xK#������$T-�����}rB��X�2��ׅ$��9)K���6ܰ��Q�h&�M��Ǆrġ��hTl�?f���)�ė}]D)�^@�M���1)���7j
���V��̟j�[��9~�d:EL��%���nK_R ]R�[�(���e��|t��n\sX�2��hbi�s�?#4�Y^�x��	��D��  u9�ϘV�4�̗i�2��찢��u1w�#�E��G
:��j��UK�'��9f��O?{!7��#��DǠ #ʊ�F{C7����A��nH�tϾ�&�x��Ʈt.Z<1��99�1����)���e��������m�}+��0�Hk@6�d��y�6���%ty
�09���D�W�{����=���k�7�c��!�p�$��ʆ,߻@֮��e�E�,ޠX#zH��7����y�.C�b��l�YcPH*F�Du�.�f	p��h�I����=��}�)(���%��Yę����;��a���I��]�j�B����<�B�E�TDʴ�*F�:hy�����ƜS&����D��/え^��t8����1�?S�+�f^A������%j��h��߽*ى�2�����DQ0P+�َ3w��>3�um,!��F�X�C*�D��4t8z��k/)0����䎭��09+�brR[�i�M�)P�	��Ӵ��]�,�[$��Oꁹ�4�!�I{ٌ���T�Ou�y�H�t�'@m��uZ�wa�nQ�'5�L�Q�	ZfmJ�H��u��c�n3���Q�fD%͉����"��B_Q��8���C!r*kz%��Ps
������XC���ۺ����K��"M���-DԦ��'~G��'��m��r���b�O`�짽�"��>A���-dr�xx�XyG�~�f�jL��6�g��q�3t1+�-;l}&'Ãt�@�s�<�WU�HA�!�BD���v^�ɀ6�(�w��b��u�1;�G�S�1�e�*zs]*������*����Ab��W1x@�Z.��(�@��׀3؊ �M]��dh}�u�!xx�рU�đ�hGr��LW6KN{�M��u�d�7��(��I��w�����B�}�S�����YA�Tu�fͽqO��KF<T+��!$��SrM\+g�8-y�YS��$T�	Zm|�@#�7���?�i��@���ܸag0CD��z=f�(���Dțb"��y�
��g���p2����Yۧ_�/�無����J��_�?�t�֜�,�`�ܗ��(�,*�gC�?�
~�܂�H�mZ��@�I�_����uU|7:��6�K���ण��@%��1ŧ��8y}�icK���E �y�V�t�w����o��տ�$F_�7>� F&
F����I�3�}i����c%ֲ���oS3̷���n�؂�j�,�	/7d�+֑���R(Q�?�\�Pe�!k�g�+s�T�K��;��+����������
�/G��.k����UeHqR�<�|�Y��ܦ��o��{��dd�p	A��?g)��V=�##�8�B,�[���4��B>b�ŋ;��c��ӹ)Y����y8
��;EC|�����$�/����*�3�8������f\��u�:1����>���^Ũ�c��K7�|�ktN/X�(�"��0�7�BQ���>���ž�`w3* q��@���9zr{J�߰�FY�'>����z7ܖ����1��Z�z�7D�/�+x��x%��`����tN�!�<aDP��&�{���pR4�����9�B���@7U��`��p�i�Ȁ�s*Ūrԧ� ��ز������w�<�+E>/Y�
;��DO��T���\5�,V8�v���q�}��ϢB�����:�a{^�	�n��$��즽8�X�vǛ���n%���^��L��}�j;��.�cŚ3ZelQs��Ƕ��k�a�=��e�QO�f�LyJ;C魳^�"(��CRc6�lZ���C���,�k��pe��a�%�3q:B�9���߈������
�)��8Pw��*)����Y�A��z(�����4�o_�-�$�Zs	X����5��a��<Rq:����'(7��&�����'�C����;�aǅ�a��p�v�X�)�F15ÖAvAF�xY��n!>�@�s�Eܠ-���A��.H�20�w��4|G�lũ�6��i��.��4o:u5Y|�qE�n]=T�
��rˀ J��f�b�Q��re�M�D"ډ�z���/��O�.E,G�܍j�lSٽș��I�^̚Ϸv�4=���|up+^��(��M!��C��=�c��v��o�K���VV'b�ᄒ���Y���TXm߀y���Gǆ���)0��V��9x_f�ǆ+����.��$jO,����o�� P��(l�X�n���_����/E���T����dQ�k�g�,�O�߉l�����2��մ���8t鄞���8���!���+T�GP�I������8��ds���Դ��fu�Γ����f�����2'm���a�9_^���*�O�4ȣ��a�`���+���a=A���}�����كAINB�'S����*��RwP�u}O/��6�@/���=:�H������;��ݿPO���v~��Pt���l�q,K�a;�C�-XKM�O>|'�"!P����S�)� a~�G�n�[K����-����ޡb
TOf��9~Mm��5�v�V���X]�J�@P�6�b�'8��y4����eH�k4�Ih6gş��*bM;��@���VM�T��U����/�9�.W�3�B��AU
6H�{�`��MOm��{sݝ��K�D�ݢ� �!����f��^�Sz6]�ls=n$N���eB�"汜�}��krO�hO�Б��*De�ƍ����|L1ؿ�)N�E�@x��]u?1���vy����k,��߬�|W{�\�����M9�U�@�\�W�ޥ�Tu{�
S$��M��{ Not��2��U ���������x�ܺ_����P��A��8�L�ՑA�Mpݍ?��Y�"�+ޖ�Sl�C,)W����g��dWa��%\k�$O':Uxr�.'|��4�Yj�h���1w9m$�/�m�)��A7w�A>z�r��0�[^���� e�G^F���E�>Fi#�4on&���ע��y�J�3��Q�ͶfB"�D��M��2f�^1��P#��̓h��Z�K2�JW�M�|쬟�Z�96��@�HJ�AlY^E�e:���\XbI���O����ZuȤ3��2�.=�y,ϼr����0�ƶ���j�P������M�>-�+,���'��{���d��Q�\�)�qR��b���6R�L�� ��T\g����-���4�tJ"Cl���ȟʹF��K��N��k��pd��J� K��T	$y�����q�y���M��
�j�J�a��o��n=譎tոu��g,��ohGb�V��Q� �Ps50�k'Gy%S��<C�	f���L�:IL�$���i����s��)�"��K�}ԩ������Y|.m6��Vj9^`��@�id2����e���lӹ��\�ꔯ�?���8�Z��8������*TP����mi�����Hdм�x�c5�A��.�Х-K��d�����N ���!�ݮ�L;Q� ��Q�=52�8���-�` T|�b�B����+A "	��� GF�#�z3#q,NuRF����w%k��a�x��L��U�?*�������X��M�y�ְ�W����g�o�~z�]�M�3�N�uA�'�D�9�()S�/5
��z(��.�p,���v����5U�x�Ǘ�Mv0-v!�|�{h<S���%��e
��}��rj�6I|��G���e�d]6{��(עRn��"j���e����}���a1���ݷ��%���]��QFN5���ho٠��2,�e��Ft��xN�%�EI��.��6%MH�6��܎�{!xr��W\�ʼ7��	tη�g�l��௰ گ% �x�#wHp���?u�f!vp��lIClʘ.�6��|�ѵ�|��a:�F��Cj��w<6#��>n7􅱸����]@xOG9"^mt�lAa�l$�o*�����*�w�4]R��D�b���:��й�$�7�� R��C.[��9j�ͮ�o1-]��]ZA��Tj�w�+�Myd�h����'�jL�ͷ��
AK�V-&a��Q�o���FE�YpM��KIB�YQ�B+����n�QC�-��8���k#Q�Z�?����;��[�Ń!<�Z�i�	�Gќ}18n1��M^0�z�g0�2��p�B��V���P�Jf�Q~�QbJFyh_�$w��.�2��y(^-����Ω�Z�����6�[����E�"&y'�ɢ��2d��N����(�q�U���Kl���B˿>��?�"�&������6��.��n������������m?�iW�'Vw"��k���e6$�g����3�B���^����{"�\_èU�E"e5�*�[�K����bwyr���y��iT6�2bp���xc������^F;h4`�z�ɽ�"��> ����B�Rf	I�^�F����)�1fV}�:�'��s^�Z�}$1�x�r�y-�VR�Rƛ��0Y&>Oo������R��r|},R� 埪\f���Y>��<4k����}BD�0��K�HF�[��J�T��FV��t-HH�9�P�+�B+���<���j�����L�F�/eZ}�vw�n�����4�q���C���_�)x�㐪h�*Y�$;�Im��7E�6�I�dvt���K^�?œ���&�I��=Ln����8=j���:zY�P�O�$V���,m-sJA��6/W�$�")�j����ɧu|ߤ@My� P���ݡ+�S�Dr%�ݮB��4�]eћ�#,K��z(ɡ�tw�C��k�^�q�� �I��gx�;��c�ؐ�-	 i�o�2��K�_��oc["��v�������fv��nT�P3gQ���f�����9X1��uQ�hۤ4��Р��N��y7��'��7^��t��lKW��n�)�9(wr~�y����ҏ]~���]��^���V�0u��;�,��۶���S��H�(����✄췧�h�����.[K�Հ]�6����Z-�����LA?��!O$��u-�%��7���	sz��c�`�2	G��v.Q%���iݳ��q�p������"rP�e��A�<�>���[LK���	��ӌ |ʃ�>,�*C���<�B�N����/d�*�dX�vҤ	�9h�BUb�㋦
A��n��AFK��l$�%����{�SV;�c�؞s�b�e��Z���?�"�_? �����6��%v-Gb٬ �9p�il�{��2�M�ױ+[�yM$�
ߨ ���;�O�,O'��\`�� V!!��&��Aݧ-ĝ�Q�b��<�uަ�n�G�UЪ�2��>� ���ǂY˵/�2B�,�^�\�6�]�E0���ԊR@�i6��q.e��u_�����;��j��o�'~t#�dLS���i�|��g�Y���A,�0��p髩��`�A�(�8*�|���| �:4d8�c0%-��	���&O���Y����:�E̴��5�qO�[P�g��y(�ǿ�����%�Ɋ��0{l�xϭDLx��V9G�rF5�c�������f�B���!L��F[e��R=�wN�K7 .�`��ľ��Tu��0K&�P��4 n,���5S,�=,m��<�(�e #�8��X����=���,�R(��������}� D�].��##i�=�g��1[�)�!&h�p<����Er-C��X���02�7�����,��w��H��14�*�K�㩛AB.5"D?(��e3F��4iaXM��;�
����)a�I�e^��[�8�Ǯ�C���RM�y��O^ę^�������"@^D�7�1k�0�R��\g@��m�\��ٞ�H���U�Z���"���%	��Q�G�����J.��M"4�{#�=����t��  �a��7�\m�5v�iy�ە�ȀxJ���>���@DɔSu��� ��&�0W��Ko��4K�D�Ұ!������d�u��5T�x�u��}��K��B�cp9B�)ǍR#&�C����\�y~�t���(6�"�r.�78t���T\:�K�}P���E~{%B:W�xH�[)���޽5!�O]�����r�$|G�<��u�x\h�i���;fʆ�����XK�&��l;�ތ�P� ��� 1�s:����B��$$t�oe�*C��4Kw@opm���Sn�on��c����P�^�d�8��͋��!}�K/;*hg�b�$��]n���a�+�����ܣMY�"0Lj{e��P������@��`3�+�>bd�'z�
���ײz� �����2��Iz9�6�w+"ܼ*P�%�d�>@��O�|�.9�_���˜h��B�9��~ګ�F�X� *:�)x�F}gLk�(G#�b��Z5���(�Q��J���o��v�JS������?)�Y{�h/�Ց,��C�r��]=���;jC�����Q��I��8�F����d0�,�V1[�߸H��Fc���Y���G�#��u�ʒT�#"_Ik���󯸡K/qM�*Ҋ�T��OU?��+�-�,|��P OOF4]rT��ܒǄXѻD���������Ybb܍�������-��޿~@�a)�;D�SY!�{�&�K$�'Y��@���:������,CL��Z��PYͷ����s��j�NÈؽ�a�̟��3Z�f �v0)m^\�R⼊�0 m�m����"�9DK�3���t(�{���*7���d�����T�4V�f��>��&�J�q���J��\%�bl�wq��G1m7�.ٗ�.�v��j!�R�DN(����+�P������E��3>�0܅r��tl-b���q��&�����l7
���0� ��	���n	���L�,��W���+���}$ ͫ)p,Py��IT��EZ}�39R�~�G��/�3'����_���K�8���z����-�����07��Z����Ff��	ex8L����Wk����0���{xȇ`*�+������{Sj�H$ABW�WWQ)�6׍mI���7��h�:.�?A�K�����É�6��������e�<6>�V1���{��`�u�~������BF{q\|$+�Q$��* �`K���SY�s���XKN��x< ��R����t�[N���� ��3	}�H�T��n�W_G�O�(lkL�?u?e��o#�b)�xմ ���^��fF�?ʹ�(G�.�/����mȍ/�a���hBii�Z�%}EET��y&�����whř��&2��8��S��L�Ol#�a�������@�8�/��;2�<S�l��H��xAkfH�_�����?5]r���\?��QQP��H�,)�%5��Q-+ף�RQ�j�6�ə��!?���1uP���O�H6�A�_�+O�2C�-X	]�BA+��b�tʥ@��;:��HJ��'z�����s��F����=�5@h���fh��8(�w�zs~� ��#~��ه���6������i=n��۷�.����s���&�bx����o^D������+qmE����0kd�o�����*P�/}�����˒�W�?�0U%���LmB��swm����XP�Dt-�8�\m{��W�|/v0C�J��ϳ��_��ꍀ��T�c�?Ƌ�}9W� d{w�n��Ͽ�2<F��LٚDj#��(��!�[�&�t�յ�K� u����~��dL����!�>����0.���+ē��G�.�bZys�b��'pZc�������F��S��ݫB��e��u��sCTܪB��˯T4�b�U�1�qf9�U���5���ݪ�߅dȒ9w
����:��l4��V��U��D���4��
E�'��#Wm��(��2vDTa�Q�rr�t��=l 6 ����I�� �6F+ؿl^�/*gk�����{gL����Ϸ��5$9���仯e�O���/�r�&&ФÓ��\���]N7�-)�?ѷ���g5iV��3G��ՋZ��N��S��3����L!����^���$��t�U�������~SƾM�9�m����+�ɐ��RJ*�=\���~�L	+����X�#���R�k�������P����Ħe���忯e��m�q�rp�>ݕ�Kd^\�1Ut�?�y���)����p	1V�Ļ ���5L7�g�[����t<j��3C��2�a1m�]b��¦���)q9QcL��6Ӓ?�[c�_�Z�\���������2�A*	|��xu_d�Wyr�N�r��l,��VME�c���44�
��o*&����)A��'\�i��^��\�d����,RJ��Hٷb�&qbt��we*p݅�@1�'ԶԔ���1�t���}���M0Pm�*yQ�7�Ҋi��8��
�5�s.�k
����ee	Λ�b|�S��Zc��R�'$�9��Z�3�]]�݉ ��lH#qg�&+�G��tO��H�*�q��e��6�3��d�m��&�EF̓�� ���^�����7��#�f8P�qp�� Hi{K�_ŉJ�D��w��,`)��h��\�t�a�� *��#�*�X�~0����]���ƛSK�#j��Rf*�0�	Ng�==�D���9�$��h��ꨍ�f��Y���L�8��t�Nv]�OU�˃�A/.(�0���2�������5ԯ6�`�����=Һ.�`@�sD��q+�^��Sow�z��)���Ê�����\jT섕���(���B�"UU���&U�F�0|���
�]b)�TB;?��N����;�ũ�	t6���(8��#l$f��\k��ՠj�3CX�X����*W=f�'�)��D��B�RA�E��M��+� ��?�<߭5�ʦ93��o���k=�Xu��N�΁���ޘɉԶ�d��5W�t�? k�w���
��BƝ0CT���MT�8u��sG44'���T�m�J��p�KE�i��ɪ�G�p@W�K>6�76������7y�V���ƥY/Hh������ MPx�j۱2���u��G�b�sP���cj�`�����JD��ҴcDTZ俩�+::��c=��nDY�l��^�O$����p��D��	r�r��`x���Ӎ�ۤ Z�K�I90c�Py�!ͨ:(�5�q�l~T�:ɕ�*�� A"�	%,R�na������@P�k>��Wj�A���4��ou�t���d8!<v{�����'w�6��cM\��_�m�2Yd7g��"���a�;󵞒v2�M �f�;?���c��`w��*�Я�0z�y!��Qj�u�Ń#�0��0��+����d��,��`�����}t�[�Yg�)�����W�G��o)���J'>z�"h�����״4����U��Z��g�X�%���?���TІ�����˯r��j-K�z@�^哕-��3���Ðֽ�B����س�����
�v���e	Y:�\��/3�$T�n0�\t�0���qi��I0�}�@!`����YZ�Z��W�1��)�D�~�*����Rꮅ���bH���nQw7��?�Q�x���M�W,n�Y�[`Er2�����ݼ���F�`�����O{��4M?�������u�uO��,a*/���`e��×G�\��D0٣��?|%7ĸ������Ԟ7H����7C?;Y�?���e�T�� cD<FM�ڒ�f�6���Rp%!�m�B#����W�����i�"����4�F����Kj/�P.�q�l��1��-&<�N,Ĩ��Ʌ`�zoyW��
��zW������G���:���n
�L0���͛ˬ��L�Q�c�P���X�*um�d���Me�A�h���K�}`�G40rS�O��L`����n϶i�	��>R�	i�%d���u�6������y2]=��I�:�زV6*������.5�����o9,H�;u��Z��&��K��V��Cv� K�&�օN,�m[r����{�*��b�5>����i `HsL�N�g�{	3̞�$*3�gp�g�E��:�@���;AK5|f�{��kK��Iv���/���=�h�j ���Bϻe��Z�z����⿐�@'��׉�%}�&���qCS诓h:�����?����|RG�?-���c��d_�T2R�FɶL��w��p�`��f6u�^H�^ANv(��c�G<A_w��2�������\S������l�{���P�cv��6��Db����i"j����V�XBff2a.xպ$B��;��%"���c�k,6.|4r��k��;:�6��m$�H� x��@�t�_<[Ƅx.�����,�ia��G܈�R��@~���"K�#!���:ru�Il�Q�=G�%(��=���/8Q�����;&�7%Vf5�F��.t��3
*�E��M^��7=��&��c}b>�u�a󋐒�∀��֗7�nax,���^�f\%��@좉o�ʥ�R���6�u�lρb7c!���m���������/]ÌB�o>P�߫'��la����V��au�����![q�m�hB��C����͋H-�L�&�{�=��
~��I4�]���n��c���V���3L�))M���@������{�9���Z��Lk�>�c=<��Ǝ��p���N0=;��&��@9��t��_�b�<�[W�ޚM05����jC�wh@W2����+72{�5�&Ԃ������w�'d�����c�x]^3��Pj�'�@ڕ�y�CʠN���Z@�Q, ���kS�?8�3�(tI��.)Z���ru�Y�*�s��]7�D2,�}��EHzkY����@n�4n�\*�G��'Y�DD@c�E#�é�X����*��M���x�Fty�D�(ѝ"Y���d���7�qw[n_�"W���̋�<*�#�h��l��D�'�d���H��4�l�}o-2ܨ_뜲;�� e0��y+�:��1��R�qT_wo��T��:�B�(�C�d
�O��K�g�sj+��h�VC�*#��x���U��V��h<��O�z]�H����Q�fH�g�r=�����K���?�%Jm���d�T�H����Z`�?C��F���yw/A^W��N�>��7���s*'ԅ�P'P����e?볥����Q"��b?h���O��S�X�����ڂ�㍖J���ۃ���h�]oG
^�PLK'��ĖBi2�D��5BP����D�a�-�A���t��m�)+�=i��@7�]y�c�b�jQ� �ڿ��j6F�[�lc]~Ɏ�|� ��':��G�����O���W������u)���rJJE�۱��I�-��~t�ܵ�����|lHp��� j��:��^��
9MV�"��{��]A�Ҥk�ݨ�`֝2z�0�Ƨ?�ZB�xH����ZWJ�ޗ���	����j����M��wߧj@��G~����/��P���#p�͕���1j�����']�m+�Ϡ�x��-^�{����O�.v�����H���ѻ+��@{�`:fͽ�_��|�M�׭%��p<�	���"�4�
��Ă)��'<�w���t���7P��g�����jc]39l�Y��3��)����f�Z�2j�<�����!)[��Xۨ��x�ӊ�`�NS��� �s{�4�����6}]�Y�ꆀZ��М�UEz�POd�qS���b�^��w;e泥#uD���{lh�c�qDrz�ݔ+ ��ű�ׯ�rj��R��\��.4֜7m� �ӟ���:h�W���X��r�����9��ʓ���aa;X��`+s��F��eH�U��.������p`�Ȧ��	Dp�b^~\[J�n9V���~�=�t$V���Ь�­���Cb��?2�5�(]
�sa�?\Pg��uq��&���0��e��#A$%
[$`SG��=��oR|� �s�E�W�O90R�ސ2�����r����
{�e�l�*���I��X�h��n���!�\,�T��� �9$2�;G�2>U���.*=p��bh�<x�ž~�&%�4p��ZnD�H��}鲜C��k����TPr��'��w;Ag F�Uzq{+-4,�ж2T�/�W��h�Wt1M4�嗧3�[��Do�Q}�CC2Rˏ�{q1DI�j���VO
�8�ޖ]nB׷��a�y�~���["�&� $��	�4�kIPh�z��oqٔ� �Z��Ea�r��sٳP38��xTTB�鼪�t�`o���NHi��C���I�����*����ϳ�X8A�LP6���KA��Ώ ���ބJ�y�t�w^D]偿�T~���N�6գh4ʍ�r�3����d#_��u?K�E�!�lc����[I�ƖBb�rg�ޮ��a<-F���jg)�Q�6��d����~��s���M�j#(�ی�
 �{�ʴ�z�5�O�#�!�����1�O�$�@�Q�էX��&��!�$�%:���R]@�Ѷ~e���#.3�݆�D*���W�8�3����k�79e�׫GhX�<?`��_k�ɢ�t�8l`<)o�� RxR�h]g�Ud�$,�:^��5��ڜg�{�����y��a�ߺB��&)�K��Ce�|2� T��a���B`�`�=����	�k]��I�È��jg`�~�?��_l<	X./a�@ƙ㠠�|�Y���ޜ�a=7=q!r��}{��K:6�წ�Jy��d���}u�񝶑Śp؈F��C�MQ��	gq
V��D?X��|fU��:!�u9�#����g����5'��`��qJUZT[�*��7�.�4�t���U��+�3�mܡ�2R.�E�܇�r�B�m����M�lY�4�:U�w�Rf n�c7��}RsX:-2p�=U��o��3�]�$�s��cCU�{z+a�,�����q� ��L�{મhh��7��Z�#I���?�qg �]�A��48�dh��z��|����@{h�3�b�ز�f$�q3�F���0(�EP=��%�b6O�~����7!%6�3���m�m��S��6�� j ����]6���w	՘˂�P?9'>�I�96�MC�գf1ۀ�:)�؏�qэ��;<1�5Og�,��^@ �839�]�TY��48������������*�o�w� �����]���ZP�n`i;㣣҅l�}vJ��i;�;ͥ�|wp�RQ=l��"g�r鐔�%䰆'S.���e�h]�UG��<Z�䲄Jm��/�~��~苼&n�6��ya�k���#qU��b�H�H��	��#.�e8�Y޸^�������y��9Bl>���-��	:�y(�cZ��~+lq�3Y�w�D��&D�%�4�Ϭ�Iut���Rj����Z$eZ����0�?F7� ���:�	��@+�ܤ�@i�n]~I��%<$8jՓ��8��JӘ�C������h��#͊���9A���f��{�����ǫ�!pxql�rA�7O��]��V��G�h*h��(��Q�x	9�4&�xL#xݮ�/�Q:)vҧ��ԷQ���U�()�l'b;0;�f�@��=�U��]��b�I��n��,��5V��B�B�^���f����E���*u�����nh�V��PpX!���mg�#g�y��;�P��(.��o���.:5G��_�q��Ƃ��1�@p�i	0�Ê����ș�rd����1�h�G(^�J�m4�T��U�<S5�Ė���5�,"hy��]�f
�9u�����.&�㦡�_.���Dzs�r� a�y����R���.m��Xr`�k�X�fk�ʝՉ���]��J	� �V�/��-��5�Ƈ⌗�^��B~O�uԵADXʴ���-�q���*ښ�����L��|2�����{�"�� w{_7��]�#ɦ�{�
7t,N�aa��bGo���۶�B~ʬQYy�i]ze��0�GE�YCI�EC�0��O�Y� �{Pt�69���T�R3�ViGV`��c'��R�� ���K��ֿ59d:����*S�5���O���T�}����'��L=�4橼����qj8|!�$9�x&4�x��9\��m�8.{���J�c�_��R��r����HF"zB��ebDbC^Ĺ�(Q�W[.�_��e{x�\'c��<0 �0�/�l�)�S���WL��s2���E�%����u������gUl�7[�i��n��ލ���*Z���j{�ݹVY�Q5=K�D���(�搵�;Ӫ�q,x �3�S S&����F���y�fRM���������e�:?�~�v	�'��t&x���i�4�hirG#:�O��9X���S`Ѷ�O[95Rn�t���Լ{�\���T�Q6:���Y:���]q���{'�
�e��g	S��U��{r�#������]�,�Kj�����ݺȧ�6#]�B\��s������ަk��O������c��E�|��0�-b�8� M�x��r�֒�R@�c�p�K7�G�+�f�[��t$V�L�������'��`/�ß�ٶ���:��*K�G_��2���w�?��E��[���L[L��,���T��x���kHX�f�����)r���܇APh<�\�5���?���jè���z���1� J1l|�`��(�q2�i���%/W]��h="���6�)�����M�&CT��OΨd̩C1��-"+�JL��킼(�~�{ɛI�}���n-?��*~(���#�%�,�]�g1��C���6� �9Qgo���Ն
9�JR�n��A�?�/�'�$�7���(,;�A�Ne)-���zdB����d/�m���杶��A�[X�
�����iY��(	;K���J�
�A�%� Y��f��Iaņ��^�Wu�p�{Oo��@��ũG?Lɇ�"0i�
�a�E��q���/L(�k��������F� �"���ξ�~iC���r�ÃPN<�Ҹ��#���}]��-��K.
]w]�B����U�4B����=�縃ew�}kK �z�a��E
�p�6h�����A�x��W�$�z�����-�'J��{����u�'!�8��5�a�E"H��5L�:ǐ���}&�a�		�;��M$^v�]�z�⠑k�D�)�3�����4Rb���v_InXW�o�K�S�.��Ң��_O8��V�<ԹX�� ���m/�Q���-�4VC��8�3��^�%̜�!��m�xh��ȑ�ءPF��oi� EO�S��SC��]A{�IF�U��h�G�\�����v�})7{)�(m���pD�f��b�7(�.�<��e�׻v��{wlz�j�8{^�"�˭~�ܱ�U�锝z��b��Uĉ'����12�;2X���ߓ�p�I��|!e 	�un:�"��9��@9 �Dt�c�Q�}������F��ͤW��􀼢%�G a���kL���G*�9�G�*�t���9� �; ���
р0���S��+�f�T�?[��g�k2x��\Q[�?;�b���T	�DNb��קey��%>����
2�Y�1ď<�����C~�o�X!6�~��H����МA\?�O��m�������H�`C�'�xA�Y���Y�/~�S��Iu�S�ذm��F��$M����xl{k��zK9p���s����!�q����,SR�}-�a�ě����r��{�O�O�8��P��v���<�ya��p_���N#'O;/���Mĉ��a8(6wU��v�BTz�Vu��
6��.�+��*Fg3��1U�-�� �
N�Z�����h/�-l���O>�_�n9W�~O�2T?΢��u*�r1\�	!D��B�u�#8Q.e�I��)��Ͷᓣ�
��{CZv��ĺ7����4+E�*����"����s:�By��P��Q̼t,h	sQih�&%�]3r
2N�K�=k���)�n)��E|A�쐽���Ab��m<S�!%���4���Q���_�@ja�1��K�/�,L��?f��I�8����=N��&��y�s�Ve���������ձ+��ho#�)V�V��Mr[ސ�2��1��:�z��<Qf��R�8�[.���e���Ă��X���Afs��f?�'�5���p�^|>�T�;�#�� �^�,+�9�d�s�I��A�ۇ�1��k+���ձk�G��d%_�M��i��2�	��<�̿���%(F=$�S���IiNJzq-�t(���(�v��Ċ��&�ٺ@���z\�<
+V�!JT��裧��m��n���ߠB!������f������6;�P��늅�J��~��K?�V�V���q�%6�H�H���g�Eg߱�.�-�����Y�V[F\�P�Ho�D�"��'f�Fc\�[NE -M�b�5�Wh�H�N���⯋AN�E}��ސ<��x����uw������/�a)%pď���L�eH��I�oq��4�ϣѪ�q�܅_�����+H,������K��F��n��6,03����Rx�e2)�cc�& �b�;Ē��]��c_�!-^����v�;��2�[o�� u/����1�n��kQ ꠙx8�ФI�y�ɫ����H���5�oA��4�}�ޣt�O��K�����GV�.�����h�㣖�g$�5�R��H�lk��T0Bv��2��B���&3%����-�>ڒ�\n������4���f<2/
����B�ܮ���I�2
l�H�ՏA�d͏G��n���<�R�
4���;� �jƃ�a]�Y�$�=��z�4׈��r�F�$7���6��4�ݔ;��f�ezN ��*k���-,@��tO�Ky+�)�>z]U�^(�ޘ�5��-;qǉw����GL^x7e��C郞��%�G��:@Z�}`�IPd���� $x�|�]Md���/Z�K!"Ħ2������gɘ�"���ⷽ���o@�=�+�F��n�SpVǫݺa� �x�6o�64�B;�%��f��/'4p2�!#�?��������Ds��u[��A'��Q[Yӱpݎ����G�eu�����`���m��i5��"�QϖB��/oKf�����G@� ��v3�7jB ������3_�T1�x2X�`���Dv��y�+������۽���.���=	]�M�׹�H�y���DI��P�3I���W���h��-F.��(�w�(/k.�)���ɐ�J@����"<ʂdy����^L}�M���XTM�[�|�6�8g�T������
���eCC�bE!��`�ڠ���+`D5�A�+���=� @i��X��D'���X�(�� 3��NE;B_��T��K+�W5��b�J�t���	�8�E�j_�^Br5�m&[%(ԁt'�J�ߴ��D�A�_���b�H'X���?7��S{������}�}�����q���'>������eN�ez���Tv@��"��Z�k��k�9宿�Ե$&���b4����Q��ʝ	�����pmH����~O�#��	�n���(�j�ќe���> 	�]�Ce̲��-H�~���-��Wx�靧�n �4/꜇�ݫr�BTG�ٝ+�A��u�W#n��M�<���YD[8�6����iJ�`�m��.��Ѫ���ξ�h�D��Kq����b�0x�R<�O�G�{3����ۭD�NS�����|��g��X�3��zL՝��H/��g��������|D*�\3Z�́K5�?�Z5h�~'蒥��y��l����
<���?_Ι��y8hu�����䄴���`V%�b;y��z����
ݽ�ﴹ(����6B��
�]��r��T�Ø	��6���8�6�d+�{Է:5
F��8em�:�	|޾�Ӷ�M����B��D�#�RG%b�Ώ_��h����Q�r�0�l��f� 5H(HΈͩ���u1�/Y�a�0��X*[�����,�+�
:�ob"�3y�-o�ыJ)�kLĦXg��qHmW�Oe@�ޞ1<�.�M��yOy[�%',{��h�5O�.�Ը?�-&�q��Ԫ���D�;�=�u"��iT��;����~��4HU
@��C>(2��p�O�@7^��z:/���L��%����=��@\�����R���g7�0:�X��t�J��m���E�b�Z0�IKQ1��vx����K� �j�f�t!��9?�1�
�̯8e�J܉��V���"����X�5o�I�{#�yhe6Y�a0��\��`4�:��� DK3X��pA\v�2��;VuU�ͼ�5� >VDq�<�\yW�g3��0�F^�Q�ο��,%�(+�s�~�@�d�m�
��dBd��Z�7�B	h���������5a����$M�^��,䊨ɽ��CՅ7�'w��E�-r�����l��;�I�ݣ=��ԛd,U
q�܅��?�|ZjQ�r�:�|*��?��}�� ���?Ԇ�]��\�	��W�@����-K��֮9w��df�v��,��(B?﨩����GưL�E(V��xg��m��*x���i�!��Z*������^�V��`�����#Jm+�<��	O�y�dV��]z5ZY��l+��{ ��d�>ȗe����'���6;>�* B�IF�M��	�����C���-�Zwd*��]v;,<���ֲb�� Q��X!��ub��<_�m��J���U���pq��9x�ʥ��@-���u�K_f�F>�F�eB>����Cp@Bʏǌ}�<�O�>��-�O7:�RA�/ȣ�\��^�i�(&O��J=6r[�#5in=q1q���=-Ê����)4��%32��b
@G��^/�@�<���.8V��xy��������#�g��Fz������|%�]�{��%�#k�d�cD	���^tr�U@�bϓ�,H��g~����U��Ț��R���������k��B&r_�H��ƴ�����ƨ$������15�W%!��� �s(��C��|]Ks��)[��|�3��-�	�3QMHb��&�HIb�/���;�=��o��~@`��;-io��rꭇ:��3�X��[Ԛ�m�T�-�)tG-�~W�MQ~7������Z��2Aă��xA%&��A���C����p�%#�K����H����	��&\��KAc�r�2�A�%���'�Q�h�L��ۀ�u��y�u���$p	�3��o����(Ԡ�Tz��K]��i;�Ō�QY��9�Xǜg)����L�q7��B�O~�l�ޓ�Aۏ���dM��H�L���t����4���v$\��*W�2�_af�#O`�����)�ۚ�A�x�e�k@���8�Z;����z�0;ۊ[P��q����c�(�U�����C�w"�<U��9�y�[����}�U��|[�������g:6�53T�%�=yGF�[��}҃���!:�X���R���0�@gp�h|�T�/����Iw�Oe$Ȧ�g����	.���gI6<��xx��V��`sf&�:���o��� ��y�
��[�R�WfLPڣ�H���RF���Ƹ���4�����J�rVn����C���v��YB����p�t�ּ4#h(.k�уn��7*]{�����7.��C g�����re��"���)g;,�C��/Dԕ�/gAC0n$us���ꕸ�d�G�X�M�\��6\Q�{6u�����s�=nxx�����#&��"�~�{��D������W�n�{N4�/���+�����M�-@�?�HN�v�����d*�x��A@*�
�aEb�<���PV�<i���9��_		!} ��U;q\��Os��Ӊ�ƦQ�Z�M�	���}�7m��C@���8�Y�+0���"�e>e����S�(�Ǌ�ͷ��ߊX>&�:�sG�Qe��k9[�I�bG�1���]<T��h�n	r� JX��V�LE��������%�t���C���=��ܙ�b9���N�/�7�	� ��	�mH]�U�ƢO�qjc:�/�5L�L��+8|�%��p%@^�SՏAJT��Js��6���-og�RA�P���!!���"#�Q��}g�>��"���te���WzY����𢑶��c{n��1�� ��~!�Yu�M>����2�3�@�x��k�\�`�)��y�%Q�3
ßo��E�p�{Ǯ��̃�_�5�^?��V2U���9"5y�u㣅Ho9��>9�?�<�@�ի�8�<��M.b�
+�4%P]�E�t��s��F=Ѧ�f�F([Y� �e���nJ���栰��,�I��[�_���q���!^��RbÅ�;yg�X\��*
�ҍ�Nc�P��K�~{����2u��t]该���*�VYn�_��}�q��f`�Ѽ5&�/�_U�x��dtn�U�-�E%w�\Ĉ9I�1�@v;��@���m8��1$�`��5-�*[��{\�F��q��2M�)ZK�M8�२���I��o�����3j��.C��c��
C!<�u��#D`�$+RP@�#��)NL̃&Zʺx�Occbb�u�
6��/�3�i�э'd���E.�E�f�q��0-�������Jx6���`
~Ԡ���6��%l/F�C2b��NpW�$<T�x�I��Ik�y�����xmjrqBɴ���/ ��qu���$��xؤ�÷`v���G�q��.����V��f��U��l�L%UMy}[�"؆��o8D`�Ԃ��|���dk'��&�x[�%�c�t�L�H(�x��O�]����K"�z�i� "�4��bK����*ǵd�iF�]����f-c�}-�h$?�}�~҂ J��Z̼h��.G�֒�Xh�GJp�TY�k���9��������ZaI�p���/�������?����s[^�5�ߡ�e��5 �mm(7�)w(��e�m;�Q5��
��F��2x�<��c��%)���o�ە��_Tt�S
����~,铫��|rD�DI�<��W�g���nO#��%õ�6y�E#v9��i\��#3����rG��wXܞ\�^�嗟�˒Ne�JƂ�>�4��N���:���`�!|
���ޯ�ׅ�e�J��~U6BY���#[ �@,�aL-���J�#���Q�J���Zb�q�\�(⒀ bD��-x*,? b��~d���2��x�������!�G
�m��LXm��8�	�>%�u	9��j1c�M׎7t�G�ԺsVN?~�狃X�a^����5X�A;����ͅ�� ��1�'&��L�� ����d��3\;c=��z	�C���F&���Drgl��^�(��_k/7pl�[ѫ��:p�x�^!���Ǚ�ZW	��	��[A�&l��,J	�����!�z:�l2Иp0~��y�h����8!�
��k­S�� 	�G�tx�ܑفX,xЦ�
\?:�n�xK�����n=��3��e��^;����D��b���T�_�Q�)�#��[�A�5��4*wR"e�9�/���m��N��1��q۝C�y��~���:G#8K��cMғ�����t��r����\�>9pb�\J��DC�q򝷠ѩ~(X`���\���Z�1La��S�N�2�6[�ǫ�y�K��W|�V�m=%��}��)�8��)��Q`��%�v@���\�qՏ}�)��2�,��x��+��E�FO,�b��㠮T �*��Nr�+���eF.5=whƕ��l���e�y��Xʋ��h���Z"^_8	�H[��X�؎Ykϧ8ZE�6�4���K�mL��{�!��.����-O�t���F�����^WP6����A�z����b�r��S!�b��~P�A�vr_t��I�\C �%.A&Nh�P8�}oAZ\��[�`�j�U�ʰ@�����?���%.k�Y��EE�J+D���Ä�g0;��v�ac�ǐ1��=�-h��L0�iGC2�O[�d��ҬI���Z7v<R#n�33Qo�f�cP���գ%kn��L��]0Z�H6�x������,�#4������R2c����)�n�"l}#d��WG�J��Mg�D,��/[��L����wU���Eq�������4@;����UN!��s�[���#'���H��N�Ja���aD��]�����#,�eC��{o�f��U~O�e��\ ������n�#�P8[-t�G�R<�H2�D�u ��%���?Try���JS�b�aTMK��{m�����y=�hh���"������*#�iP��|�)�#�]=s/���f����$���Y�+L?Y��[	��m'إ|�}�UA7���OX	&���^��A�8 �5��ߜ�-!O�W���YA���@	�.�T�#��X�J�U�u5�\�ϭu�7M���7wf�ǩ/���3�3�W�X�t;,��M|�Ӵ_�ꫀ��N=F�����VD~ϟ[c\��,�UBaN���-��{LUŁ�dr��K�C�E~vF�%��г��DP�d��0�g7P3��s���P�A�D���7�i�ilvG��4��fK���?�̶�3$��T5�h�6�F��E��r��7�.�2J��YaWV��T��li��aM���������_��P)����Tm[����%��{�A�Ƅ.� �c`��[lp�t`�c6V��L�qh�	�2.x�����q�"K"�]�/�Y��<.�z���p�zs�lv]�U�_�R��i�VUAp�Q<{42�*�N���P�K�S�;��lS�|�L�����Ba����v
l�'r�@2���a��5BF�����(cUΡ��J�<���=̽Pa�R�#3n{�V+"hp�}���kʓ��ƌ�GZX�B8_L�r+׉/I}��Z�1Fi�֣�ek�B��>�����|)�%��35�Y�����i�F,\b׳���,xv�2�:"��1�ROv����8~��f[�3��e=�[�K��]�h)#~��gqw���0�zyZ�3�g#����U��l���O���.DSrS�VG����ϪE�W�LQ���*�0�(���B٩meu�Ǥ_��>?9>B����ӏ�Y�	��1�)1���]϶�\�zz,��:F�x'�F��_�EF�v� ^Y[݂�d�q�˶��Q$�'�>�H#��wK�=�"2�cKM�t1���2�V;�i���m�$p�Dqì���$��9NS�.ps�P�����P�h��Tf�!��5��J70�����7��~n��_^h�c'���Uot�tڶ�����ח$�1���� c�ݑ[{�¢��������б�yA��)]CiyA�"��L���W/�o[c
aВ�Z��acY��D��;��@�,t�[
�.kUu�i+�yU����
�+DMF����i( )���v�e�؞)����aa.ri]h[�ֹ� �o9j�|�P��"�+.i����չIQ�Խ�|._TI Q6bGJ�G��g��@U�C��j�7��e��Bŷ,��&9P��w{�w��"�>¶y},׺&����P��.!�4��{F�a������8�˨�Nc��K��/�����TtbZ�$��6�Τ�a�<<:��)Ϲ苛O��H�ez,*�>g^�J��:��f�
�*�Ow����͏U�5�2ُ7�é�H�8�5E���M=}���8XX����g�2��C�z��|9�u�/9Kp�u�L��iJ��}Qw�EB��b=��&X�>�A����"�8��P��p�U�e}����L���LQ���B��Vt�z���@���)}\��1�e9+����v����L��u	�����RxWHc��v�򌼰t-Խ-�+p�uȅԬ�V����a���6��F�{�6:�SS��Ck�q��&�meP43Yl��X^"�.����L����B��5���+?j�ե �qm��&_��M�ۭ��i���`����?*(�p�;A��bSD����Rʉ�}���dl�=.��C��&q�Y��S�2؝ĩ�K�0�= �I1|���]�LW�6.)-#av���ʪdn�!�)P#@P��?\�'B�7�DLs��8���TK}��4��b^����tRT���E�B��n�nG��&�|Pдu�h�B4�t͚����ş=���!+!03U#��-�cKب�=���*���r�K!�G�
�C�)̳l[84��6 w�V�&�E��-�抛19�KMp�����ƪ:$��h�;q���0�5_@����ܾ��C��H�cm{&͖)��j���Z��1亗�AY`�� Ł�~���q�#7*g�g��7)s�5C�,DT����d����`\��)���p1�j�tõ\����(��l
`����d������k2��wQ��C�l�u����}��R�43�Pʮ"�s�to/k
H�T��&�U�3'5P@�1=��X3� �q�%1��Y��E�Q��D��j�����Z�޼�M;�闀>�����d�s�-���^qh�h�`��9=�~�G�+��CS������w�ZX�p�c�������#͸eL��R��M:u������_���m�0��e���%Z&ڂ�5	qs��d�10����k/t�a)������������%��	��q,z4��B�HC�8ŕH[��05]�C��aH�;�d���ɧ��h��c�*� xW?�\NFU݃�I�!#�h��{�xCeT!�Au�7�}1�!�K*�]��F6t_��wہ�([2Q���.#	=���6�������2�b2�|&BsB �L��vh7T�:i�ϯ]���K�W���,/���e����F̘T��Zl&�jq��pީ�`���UY����I�>ɪ��SNC��r����$J��f#<�x_b�*�,�K��(WLXW�-<���KiL�Qʅ�]�=������Ѳ�K��J�Y�U���3��)=� 8� ��¨X�u��V���a��Ԫg5�������n���Hfo5E�/�ua �$T.E0��T���L���D<�<���&���|*���m�cc�~�i�N��2I	(���Y*&Ko�s������2��hM��G!T<�;��Zv�^���u�*agL�m��|L��v��KV`ݧ��5��"�Hֹ��a��-�	>��=�0����7���Աa@��4A;�; ~s�}�[��5�.sE��o�D
m�KuȂ�P��i��˝]&f�����xH�_�2�&q)Ov��a�p	C������S&��O����6eKb�8��ؖ�|4(a#��!����^1�.��ΰ�q��$B)9�k�m����Y���"�z�y�5�Q�}Hߋ9Ǥ��C��[&%p��)=�%Ď�W�r���V� o�F#��)�j�?�W���q�6D|�y��� C����1�-���{7W3!h�%��]�n��_�c�z��,:�oD�-:�#s���46�����&ȨF�wDn��ZD�8�F����UH�3,Ю���I}k�V�5>g��y]�ږ�E�jv�	� 	t��1f���t��O�<��
�gֿ���TBP��f�P�y_>.�F2?�!�<Au����z��F��P-�=���g�����YD?8��t�}3^stpM}ww�ns�OT���ꆷ3qBFy�cNk��+�P����#��ɷ �KTsJ~0���x73p��e���)@L���]�H��:�>Eh6S��қ�_<Ǫ�c=E]����'��$�^��C��o3i~�5˚e���#�#��jg8��A*m:'h����u.x�����E!��n	���n³N�`�������6�c��N������Z���8.F0��++	���"��������裀���`�.�;�Q�ld)DU9@�ˠ[�:N�-0��Ƃ�����YU�P�D�>��T�I �*�c>�W�I�ܻ�eS~��?5g�`�߀}q��jd#�|����V8?��|��y�vt�J<%����,^d	�[D���Gf-���5�SG�bڭ8�b�0�y�O�]'w;i�Ț�n!�J�K�oe�:@�>�c���@Ǜ�6qR�￳B�C;쭦8�\)�;�D�b����s�d�{)
Y"�>�-�����A03�3\&8���f7����8��iq/���\Sm�ыj��U��q)sq����E���Tڅh"�uw~şB�#�Y���$ՠ�_iٌ�_Ֆ/���	0("�x���f�߅�k���zZ
~�ϙ�	F'�%ڞZtGP����oAb�J�8`�D/���Ǡ�;�r�8>�ح�?t�u��q�y>�ͧ6ȺwKT
��"��Iu�f������� e}ۅ��p�L��Z$t�	��G���d
9��� �W��"�>p��b���c=]d�\�)��,$�]�6X+�~Q����65�]u�x�$�PB��N�Z�"d8�!�eMO���f���6���5��?L�*�*'ú
X�2N�:�br ����m�I�tP��� ��Og~��vQ@%�3���O��j�|\��F�b�JQQڼ�ҥ��#�T��\�I`�������:��0����I���[�M��u���_��ȥl�������Ҧ��֭��K��a�����v9K�?AH���m�(����d}�&Vu�o�TV^�	ҳ� ��ԩT\^o�]�O%��6_,y����5(2��J*�&ҟ;�
!�^�`����E48(�*��9�s3��B�������i�3��&��>���¦Ca�,�v��>?d��~�˽'׫%�{9�f�hG����H�w��~�
[�8��T�r�w8��#߻��݇��?T��o�Ѯ�ʠ���ۢXc텳�k^�b�޼r1/M0B�)�C��0F@���o������MQ9���V�Ŕ/Ծ�v#Y��nU]X�ܻ�b� �_��D�*���T�Of0��{9S�'u�ЮM�]�u(7��w#c�1@�[8�[��"�gD�}��WH�����I�������;�V��Z:iύoc�nC�i>���W���	�ˑ>���$�`��U���]]J-ڰ���7ج�JHm�Y�+BË`=t��My�B�
��J�St�-�$��|g'eͽ^3�
o�a�=p���j��_ݓ�h�'�r�j�Z"ɿ�Q����x�ݬ��]�G��`o��@_(�^*���z��hiK�Z�h�U��M�Zڳ|������}Jӹ'�q˸s٦H\/���h��](�	�uK����BS���˪���h�S`�1�������9���1qj+.j��\��i�QEp�u�G����^�����!"�8� ��i�#W�P&��F��E��x�=⅕�<~����Hdh�F��8��l����(݉���*�&s*��2g�Hu��}7m������b6�}��򒢏Z�vQ��B�0��Gl�j��&y��6G��$�d����$$Tl����P�i�������O���ה�zK�Q{�A�&�<K2uC�mхx���@k������ #�IZ���m�gH���z��-���g?�.Z}�c�z� �?�I"HOG��>�8�ST7�9�%�Ʊ~dl�U�*�jM�G$S*���qߓ��Z�n���O1C��3{f�$�'pwH-��� � ��PoI�^>���
�ع�=�W2��u�}���[.��0JR�n\P���c�$Ӧ�7�&� R]MƁ�L*��{S����02oT��_{}�O�|芗&̓��k��.�q����L��x�*,h�P��:a�}%N��}p�����l���#�u~��H0P�8ȬF4l0�b_��F
��Zz;)�`��g�x��o� A�x���w=��Y�	���laS8�J?��WT���l|�z"hdHCa�V�{��A�8�zה��N_j��J_�5�CP�M�H$`>Zyc�K4�ĵ8�J��a��~��W�K�����_?1�LK���������*.�X)��`h�}yݜf��_���g��'��˰D�)�����g�Heg���+�ϫ������+>Ҹԍ��!
$U3(웪��Ab��:�6I�U�lЏ�����Rr��u���'�,����W{^S�����>������뜸�`�	�g��=)XU��`�ܽ:�S�Y���oi>u����zg��1����~;�WFw��
Ǳ��A&����ϋ�1?�9VM�.�"D/����'@ f<l�?��we>"ZyL��F��_qS�6T�qPA��)F�Y���i���ן�UD�v6�?ܗ���)�q��0�v�/��@E9�X�0��8:��D��/��?��@��-"M�K3Ǫ�:p�_�3>-9M4����S�x�'�$Gv�$����*�^��-��*�-��5�___�A�-��]�V��U���o��|���y��E'�请6�-J��N��%W�t�Xhv�ذ҇��ˋ'^-�V9eRk7�2��15�����V4;�&�� �F(y�V�a��l BaDd=G�l2��-����#�C��ϡ���"%^�ٱ'3kY��/�\�w�\tt^�	������S�Yd��%�Vӌun7nf�s-Sv��=�;���B���,CHJ�fԏ����>��ՙ��ʛ�>��H]]:'o��������ɪ��R��ҭ�����t�p�5���]D�!�A�6��]����:x�%��#�x4��61��$]�*�^;�-���wl���	�jo`%�l<5U\�4�;���x�3��e����^U���P��J0��c�Y�/2���o`�MN�S}�_���*�o�]6�� ]@Q;��l͵�f�rOѭ�4���{�ʂ5�|P��D aH8�.Ր���c�߂r�Et�I�L�ӽ4�������S\Y���B\���[k��⿥O3�����#�@�X�	��E�X܀�)��ѠfE���zw�ڍ�\dU95	�6�D�PfǑC�� <��Q���E������,Y���)��&F����<<�O����������X���^D�Â�d��"�W���BxH!\�3ѿ��W�~S&����qa��>-pyzhGS�� ��Z�r��lD\�.�%�M�Q�T��=���z�'!��J���M	�4mT�^0I��aaZ0��(��4��w����Q�F�H�xq��Y
�wup��mM/!����UBJE.J5�g�\�pX2>4/��.���fK�l��PB���}�=M(*��2��k�w�p*	,��f���X  ��@U���f�q��$���5� ����'׌ͪ/�[ ��um�N��կJ���#Oq;�q?[�!��ו��c�1�l���9ʚ�o|��d%q��M*\�d����i�6o�d?�f[B��$���?�ƞ�]���O��6�$�s
�?c�//=B�l'���-=�X�Y1ͷj!�]�)u#D���\�2 ��|>�h]�&��c2�®�Z���~Y�Cp����8�q=���(��N�~٨n�T����%�A����F�m�0s�\��d��t�^v��rڵ���c78�U#��8P|
+%$<�ןЦ]=��`Q����.z*���c������n�G{�n&�����!��]�UA����wY'ݏz)۶p�T��)L��.k&� ��/�â�M��y�_�P�L&äeu�i`�t����b,�$�t�u�&
p�4�65��ڍJa��`�އ��I+��+o��#(c_�ϸ:r���s��e��F�J�X�}4�����|�wX�0/��������U� �ҥ9BG�Q- �&���b��`*���S[���NVCp��玧#�I}Q���U
WD���~�+]�IE���>�iP�� J@�b%�TF�Q[���q�{�AC�?��4��=[�mHT��"�C)\A�����cCq��S�Օ<�Om,(�#�7�'��^�\"����������l�ʰ�jwF'�W�B5^  ��loIkr��d'��G�r�w%S�6��B~N$��bʓ%����+H����nS_;��M'��Tǻ��$�.U�5}X~��c���"��wT\{�<|+����h�"�/�,��c1�S[�0��+�GO�k�Q�LbWO#��˺K�H"t�f�*ɩR���2��W�Iؙʉ�M�Bv�j6>���7���a�X{���9�N�m&[v�L�8V��^��]�:>��wy�;��SZ��:>�}4�:/��N�!l��p���ؔocC��T����^��`��p!i���i��\/:ڷ�\Y@B����3�w���(�#b&��_�g�uymz��c���Ԇy8b�k�x��;�(��g��Jyb�,wK8z'�M�$B�*���ue�6���p/�E�<�u���������h}5#2_����v� � �{؃M����H����V����ި-����m;;�[r�WM�^�@㋥Fۀ.��h����g9>�����R�H>1i�h��伜�OD���zE��J����M�!RIB����JI�F����%�X�#&��^"3�9���W���*���]�/���y]t>`����ӱ����	M����^z2I�~�r{�����pzt��s*hX��/R�`�s���q�t�P��*fz���X�f��>bx�p����0� 9�{Mf%��Bם��u!TE������Jw�lؗ
N��F��Bb���)M!�m�ﵹ!�{��Ȑ�<���ߺ�TX����`l��%[�e�z�Һ�3�3���['��m2���@����`�o����ݬ���逑�L�R��"�V��b��o�G�h�V89p�z#��h�mg8�ұ��7�iu�אx���O:Lm��`/F�%ms�@�1x���3[㍯�c����[S)*��&���S�#�Uk|�37�hA�����d���w�� �&`��ֿ�L/ґ	|�T+h���P�R�Pgz0���KK0f�w,��k&����Vyay�Rq�S����d���/�4�*(�u��������NQT�%��6k'n���:���q�����]�
!D�e�ӭ����z	�`SQ�U����H7�V\��ߖ_�>����+/n�_ S � f�u���eizuЬ����Z°s��#�΅���ԧ"P�QDR��΂����3��=��z:�o���V��ol.�%����4�����9�)=Us&T�4Ji&ݐT�őwVҸ�Xҹ��{a�TdC�I�)�Z��\ w����ʙ��xn$��/c�if�H��	3���Rg���9��j��њ#�c!~�kw�܌�BIݡ�v���ךI��>w��@:P�¼�+M����T�c�⡷YWq��E������ކY7*S�;m�������ߜ�ȶ|�N�Qz�^(9�/O)���27��J��*��/3O?����y�����Q,��&�t�O�G}�9���}r�U~%�,5,�N�N�@�}N:(�� P'�@�yrn��|FNºu�l�]��4��O����80<��y��
���E�s�1G�i���N��O2���3[��KL,�p����e��`P���1�w�<w��t�9Wt@�q�tZ��?���Y���zld?[S�� �t�Ql�moj�F7���:����)��Ӎ�\(h�o����M��3єr��NjT[��G��3S�}���͙��mPe�5�$������e�5Cx����� ��?�1�k����)������bHվ���\�WyL�'X����\A�A���\�Q��1 >����PB��@�$�B%)W��L��r,JՍ�E1V?R��U#�6�����GW�F#80��S韌�A?��u�\(��^�������F|�6B�X}�(��6�8��?jQ6��`����z�]�4	>K��,\l%uw؂\N���q�<a.X.)ܕo3�&�e5���ߪ{��"k��;C��n�g��y��$!���s:?y�2,F���VC1��&#$y�l?3U��Ҿ;�}�z��
&�+�Y�:`�hz8����2\��cO�a�jw`D
$�\�\p�3R�y�.�o�V���L>��+v����N�z����`��s�����Se�G��l̓Y�7�?�&��<��B���U���?,�],��払��٨H�m�y p��o+�kP)��S4��+�1;�pXE�I���4q�ԛ�d������i���	���e�����\����;��?I�MHٹ��[�ǅ�%�Y��v�LdN�X�A��H�[�m<��H��x���9�4@�-�PS\��ךlî͈�nhh�F6fIjw^#[�6�8�WԬ�D�
9�:T�I�lg)�q!j1T�%�K(!�S������dLk9�8׌4��|inQnF�;��d�S)�u�U�w��7�����~o�vߍ���k�w��2���;}���3���5*O�>@p��$@�0��*�8�@��сV[��'�91����ȟl�:8��PtH���wt�I^X��F�}�}Y���ז��͠��'bd[�e���{��C��۷cJ.��f�Y�+�<�ޔ�1wM�� ���WzX��/�;�ry(	qp����� � /���@?#�W��;Ub�P��՗z>�36?*wJ�L�?�M[Ᾱ����nJ�S-F�z�_��s��!���,Ln8�#�u��d���4*��[g��҉� ����SS�կxi�s�"�W��h�Ƶ��9h���j�*���idQuЖ�*Y�Ը�[eM���k��6�G�p���d��݅q�o�T�C�?t�dw�#�L�و4�����7�}'Q74
�R���B����#�N~X�W#�z3���-�g��r	|�a�g��7��.����(hr��Q����R4�y<���� �vqcS�3i���"V�r�~��["=s�d�����闲nk����f^׋�ư+�"@	��mE�����ڝ"���s�Q|���)<Ԥ�1J��PsX���8@a�-��?L��T����꾭w���ރ�M~���7#a>Dx� F�H��g�Tz���겣`�n�M��(,�i�`����
d��S�hPk�TuZP�$���]�!� ��HE2%:&��v�}1K]觧UeJq	.ɝ�&6�a�[�^|5��{��O�Ƀ&���}�����tJ������@BR���cU����pM����v���g|Q���R����ʢ3%+7ѵ�5!����ܙQ[��F7��g��|T�k(�E媷f!ƴSW��7����+ez�X�u,ci��
T���i���!����΂K�p��k�e�����5��m���3kUh ��l�n��e"熥����
���o>|�� �J�$��e^�Ι*�x�����/�C�e�J����Bor�,�ҁ�#��j�r�g�Dُ�OL� ��/��S�~�I�X���� �:��ѭ���@.���)E+e/��t�]���"-���<�2�L�A�~u4��&l�l�Oo���-Z�2�F����F�)2�\�l�[q�GR���(81R��ъ�ȮG�S�cg�\kseT;�l�U�4l�P�*�P��Нq�$�6�S�˅����^�ћ2W2w��O�ZV(b��6oZ�����o\\��qp�1���4�hk}\}�?���q_!ƪ�f��yz~Z��l�(<����P��Hh5�y��wW[t��Z1-��g��HG޸�P�|%k����[�U ���[^��ʽ��F�2��lV��Wö)�
w�uN1�0�	2������=y��y4P��nDɟ^�2�vzӨ�d�	$LW��~� �X7+��2����>��aM��D�t��#in��3|�fο}���;�0�5,��G�����׈7�����B�;��5&���j���v�ٹCʈ:i��Xn������V�r(�����/޵R��c�_"N�J�Ԝ�U��T���~���@�XTB8�X*E/�y�y��?J{Ѕ1>�]�� N�(���gQ�P��e*^�8L�5�p��c�]\��P��EP
mN��5$��l	��Z��OklrMVعڌ���v�!K�� ��+���n=W��U8��b1��s�z��%�&`_��\�r9���5#?��u�Ta���g��7��V�h��rt�&�f��������H�k�k��3+����M^���B=s�2a?`4F�'��6ݱ�9c�JI���H�|�7Q��<c<*��?�`��:F	n�%��ޖ���)��t�P�I���_P���@��y�Ik����1?�@,����f܀Q[0Qx$�D�� �Lζw7L�A��	� ��(�DH���	NW�5��2��o	�k�.�{՛�ul����/<`�??��%T��� YT ��B7ʠ��O���~�:��P�g�4_��ة l��4��{���Lc�5B�;/��YaGlR�"��E�A��U`� ���l�L]���q/�D���%�މ��Q��z����,*����l"�L�e��m��@5<�e����n^�i�u9���*A�����wD�b��D�
-,PuG'(
���(��hA/C��"5��-�Z�3�qKL�<�+���>mp�9�G`�\��n��o�)v.��P2�&F�%�Uu��(˙/�9{�n)��.[����U�~`�)���, 1����%�(�Zފ�_0�5H^ �_�{N���p�C�6���A���6��������B^�]bT�-���/e�@�y���PY͸�j��>�I�*�V��ЁM�g���3PS��N'_E���<�����_���W�rH��a���@�[4��Y���hD�ux�Y�`mX4�'�Q���\����R'�%��_o�� C��M��]�����R4�pK������x��J�aE��7����qy��9dBY(*����Γ��ǉ�l[|~����,bG`����S���e���Z�Z�̦�'m$�BߦTꗁ��+K���'�Qvt��ʶWԚ�
) ���^��thHd��L%/�:Xö��u�O�3t���?e�V��$f3R������4���Π��	\� ������AVc?oc�<H����G?Df�GG /��l��?���s����U���a~Gy�A!E���n,Va�G���x2�\�;���H�ͨq��� ��BKl;%�va��#���HW�%܆���=I�{��SRfh��8���FL�DD��3���o y��.d��lE ��
�S�=�Íu�ⶡL�yӜ6��13^�����K�a����F�R�桟V���/0��.����T|����"�x�v:�7�[�1�@��`,\U ರ�W>��S,O�����pk}N�۩%�
zT>L_j�2t���R�NM���	6�v2�16���a���&CL��|{��Z��۞��U�1$[]d�B�zpba�VF�4!�fŊ�u������_?�c�1U�����H��8]?
Zu>RYN������)НkV�{�S��ex�{�Y�V��e�Io^�R-�,�<���\�?5Jh�W]�x�x�n"�&�sO	�����tun�*$l{
#��-ٽ��X3E_|�n��>Чb78�'M���"iaK�c�f\0�gi����� V��g�A�����t�Mz���f^|�PZx7�H6]���bT�����=�pV��T�S��Y��0*����b柾f��I�%�mz�

,����Kk���K[d�M>$w����,`���닒7M�U�^���5z3��h������˂wa���9E�<ϖ��w�V���F�"���܍�:gT9��sѕOՏ�ӿ�.+��;��#."^sbM���E.���FV��L'�C-Nu*��u�>�du�/��Ӗze�sX�'�� n�� ��8r��JP�U�y���־�	�UD�gy�������d�~n��K����:{5��_'5�R=�V��9�Sb�<��RIН���ru(%�>�%�5�6cKާ[Z�S���r,ҍ�0zEg6}\�.x���9�n��4�6�.e>r�*ƾ꣨X+��nH"��':8$�.�A�0L����Qw��N���u�O��W(Z��lSZ��JP��,�Mt�Վ��!<]֥1��}-�Eg"͍p%���u~�>N2�b�ib�Щ���=n����p�{a����G�  I�%��"j�	j'ufm
z[�q�̮��R�*L\�Z�qX�~Iw��/��,4m���E=�������'_���d���Ѿ���}��.>Lt�Ֆْ�7.�(��We��Ƙ��g�?d��^TA��\L��!D���|K�l��=)�g��O^�cj���#�Az::����:{�3?�8������o��ѥ�� ���\3A��RQ�@� JL��3=��a��cmI*�	@�R�>X㞚!��p/�(u9+E��(b/Kl��I�m�����FlK�$�Lm����jW���&��
6ק[ֱ!��Xd�髱���)�ݧH��A��U.�A��v�j���nj'ʅ��Cb.��Ā3�,e(�뚘�^g�+�b?�=�1�	�%w벯�ޛ��z���2�n!z��ë�w0$����$�<��i�@8�s�c�����Z���G[��)M�� Bv�b�P|ͷ��]��KI�>�`<�z/��:%oا���	\��Xz��5���_��C!Q���Kd�G=�R�^�B1u�9]c�u!���gY��N*���ћ��"v�bKi��dK�;Fug�+��"��ʘ��@��҅#W.��(-�H_����U��&�(�'��{�/>۴nZ;�1�(�F���8ᡩ�	H�����"B�Hi��R},z�|G����7�Xh�m��531��VZ�hV�'��5h�<���Y%��у�*bo�̗K��6k�j'
2{�[3'W��[�m��}ߩ�	ɏ���O���6�ɢY���?��6��[)a���4�<'� ���>�^UBgj���pO�f�`��.7a��H�|�_>IJ�w�W5��E�JՒE�����k�^:6��;9<�cw���c�[��C�H�K�TG*��	���-uk;��騼��@̑[�z{������wf7�Vc�	b4W���G�6��*��-�s7�E�0������<ur�p>E�|�#M�5���1��~4�-ww�&ފ�����GT��E����hp�����8���#ƃv�A� J8zj,�k��tI֑����Zc�����b�����'�v�}�t��v"�HO���G�#]�uOR��YB�Jt+c��,��gGQ�y��ݫ��y�l�#�ȿ�4�B^H��� ��Y�W��,�ӣ,���lKd�pq��n2%���Q��0�L�:��V��Q*Ò���^7s4�@/��b�X������9��Y�q��ԓ�d�>�L{���e�ǒZ����U �\�i�_�q!2��,����(�1&RD�%n���J�kí�'���z-E'�鬩T�˪P��1�W����m�k�c����B_Y��Y��7y<����_(�D3�%;߸A�R�z
M>c��i���mC�����yU�c�=� �@w�Yd��Y���k�X�3lhA��䨼����>�(��=��X{���զ.$���h:��\���Nۥ�މ��Z�vz���&�� �טC���Ŏ���:��e�f�A,ˆ��~���%�$�g +�p��Yg!�ꬭ���ܓ�r}㸿�r-6��t�au�Ҍ�2T�t����v���Љ(���u�P��	��\5��YaE��U˓0�KV?��7���5/,�"�:ZT�	�L�-���Q*~��5˄\�7zB�8�\�s�� �Bc�	Б.��_VF�Ż��7Rj��`�GTDz7���&��V"�y���\6�5 �:��h�~i!#[7��O�E�'L^�y !Gޞ�Z�c�IrY�f�װ�Z���2yIG`���a�����(��ؒOk;�(�a�i:
�כo�br� �.MH�*�����T��n˰��Ԭ�N=;]�1`Ŷ��Ͻ~�����l��r���f&��p7Q���*����>:J�b��y�:oivS�I7��)5T��@=H��KG'�	B�L8�2�N�u �S��f���*B��r���K)ɹ�Y����f�P���_��sU�u�Z�T,g2瑁�\y�nZP�5�?	�(ڸ������DO=%v�EG�]9"A�O�O�T��M�
��J-!<i,zL���+z��o��v���p�����+��W�v��Q��~�$�5�& �JV���-�Q?6�cߋ�X�z�
6�ɠP��I��|S*�0 T���@����|bL�̹��?N(��4 wji�a�����f:oM�֊zAw�����NѢn �v3O����5tg�#5�_<$"�h�b�Y��t�=��i\�	>+�^������R8W��k&�n��1�e.����'r��cI�μ�����6M���:E�A/�����Ihy�\�Vz����MQ7F�R\����H�$&����X�"�e��J��g�6��i
�3țc%�}%�d��NXisz'��.��b*��E9a��t;L�\�C���2��E��ҩ�r,G��bډ��=�<�gR��5_g5k�к�h�Z���Y@��KI>|�O���m��x��F�$�-xDZ$ �^I;�´U�$�Z���fx�#����M�o�c����(4|O�Q^,ެ�����2�nz*0ϵ}�:hSu3r�Һ�E%��js��4��	�{iN��&-6��� �&'4x��0���d�����۝'���i�������Go�W�|�c�!_taC_�3�l��਱��B�p`l�8k�$-���'��P�z�r���rý(K�ۼ]E� ��ږRȤ�8E��HӮ��׹�6 ���WR( ������O�.��l�P&���Q���/���ni-i�������>��ⁿc���k���T�8`��/sE�|�(��rB!)Cn�9�D ��4���*�=�3��L��_�·�e㥱!Wԟ��U�eiZL��{^ޜ}�e]d��t�h寙�\t)��T�.r���2��Xa�Ɣ��	��1S��a��OLeg|��".�3� ���j��V(v�Y���ʣ��6
��_���D���(�h���������"�6-E��R���7�v����h�����f���Nb��VD;�F�D��O,[����@�H��H�*H֣����A�
N��-��A�$d� \r�����s/�zF۷�gmh�P�ق�V�8Ԝ��_@������k=A�2<�E��Q�AB���]m�5`G�P��jU�[Q�������Q��kl��%��`�����~0W�3�0������xG�P���Y���ea�H���cP��Ž�3�WϼCbd߂� �y���Mk�':��6tq�Nb�p"^��^
�޼�{�+��<}����Sadr�5�%EA��c����8ؤpɘ���s������A�DfGt�+!��q�%����E�P�R�:tz�w��}����ڤ�[_`�Ь��vN��6<X�e�)��.i�M�.�����������<[v)pq�x!��K��EQ�{����$�u!0� ![N����6��;�X��N�Tw\%+ӊW,p�s6V�f��`�RS�~_|��Z&��߀��`�A�K�g׊|6��ʿz_�(=ꪀ��ڔ�XbK�ϜV��Z��ލ���#	��Κ�����X�^���zy5~�o�~�n�Ӈ�<�%��sw��
����V�u�c�`�6��RH0_ Ϯ�������M��>�9S�t����Ɩ�^L��չ5�/���@� -m��̃\�Rr�v
�Q�'�/h �F���y{ +��Y���[���0���bQ5�(l|;py ���Օ�ȯi̫
�/�0����"���9S)J-���_X��t����ly�F�Q�e�.'�2��[-��i����9�қ��tK$a ʈč�+v`	F_-\R>�S�d	��A?I�(8�jN_pv�Ѿ���������C")Z��R���c���yю�S_�2������f�.z1�>���f'$E-ٮ��k=�f�x�b.5'�� E��g�"v)�S��_�#�h�G����b��w#V6��ƭR��F���6��91�]���(�0��E1v� ?^qz���(!�	��7Y�p��=J}kd�:42@�n������ɦQ8�(�&��M`��N�.c|�j�z�����N'
�$��wv�GȽ���H�?RF��/G��Σ�2�>@���u��l�S[Ll_(�*3w�:uMH�l֖��p���/��I��3�t��l�~&��
���:X���R��̩W�l��7/��l�VB�� +%��H .��v8�A%�����˹�q�fȗ���T���ʪ�Ѕ5Q_J��h�3�Ek=`�(`T��C�5�g�#i����@
g��@��5� ^�QL������݈h��zs�CZ����$֮�/њ!7�Gc�Su��G��BY8@B|�W� ����?O��tA�Q���b�X�"؉�p*�\��Hޖ��Z£n ��%��5%����y�@\YA;���:}g�a�aP^5�ޓ-I���Dv�X�ܫ����g����t��f��%q��\����r���ƈ︋��j�`� ���C����ahk��7��O ��?�ɉ9��d�̟̒;��sI!5*����i���3�컓0��jhҟP^ky31�=�OKE{\��#��Q_��#I),H�:��%4���̅��XI6ݍ�$�3)'�_��]YL]�1k/����>=�V��Ke]�Q�僊3r-�Ka�k��%���﷢�QA��%��O>?Q#I������W�Ͷ���wf��N�T�/��3���mkWD����#����V��E�����68�Q<��+�=qSS9*����md���?���9a�A������e~B���Pm���*W������x`��q���֯@M���A����:Q%���끧UI�߫��HXmr�./�<�:WF����$&IJB�l>�$:{��N��H�Gi�Jn���U���^(ʕ{�/X�ۅ������R �#�)�<z�lԬ�|�lӒ�� ��(/�ف��$S~ZW�:DI
,��^�UT*j�'��#�@�8[/�eߛ��8��m=�N��%}���"�;G�G�c�h��+��U���:eR�H�+��[7
;b�c*r��S.�^ń�Ŵ�]0�<�g�3��ڧ5=x�ceDb��n{����e�)�ӝ3k�^"�	�x�D,��	�:�7�p/"P�.��z��7��!�����A�)}�Z���r3��}G�����8�d�����E���d�G6˺$���%M�K8���e�d�sRO9ܓ���������0��p��tU���Z�X���\���ʆ�+��8����m����o�7g���D����P�p�� w�ɔI�_[7*z^#�c%U�����,lᆡ}�$��zX>29��^��e�S�������4� ����}3dc����*F@߲o�����%(_ �mB� �u'�WB�������a{8o9��ta�XݥK�r���r|l�v��㡍�`���,zb)�Tֈ��%u��X�Z����P(���Ţ9�j��T�����:R�����*�ן'��w�m�#�}�Ǟ�����F�Z���DV���]^��P���Fd��Y��Ȗ�a\���Xո�/&�h��;�\f&}]�(��G���w���dȻ��!|���j?�"1^W���OSdf��q��o�:��V ߥ�;q<Ԥ����JB*��[if�鱄ϻ�f�?��CNѦ��Ǟ&��J�f��w]���$](��Ut��S�y�;��N�=�C��,�ctT��$΋�:�>���RF7���P �+��������x���Չ��T!������6�n��Y��s�2�Ve���^�b/��;��6�zz�*y>��	0rC&��P��P��d���ϖ�up Z U�\�H��%#�h��awtiJ
�c�0R�~��2y6�c֊k�	_zyt�f$&��a��$�#p~I�r�I���ݎL��Y�Z����W��`��\� �8g�s�Cɦ�'n���֠���xn�eM�������҇�!��I�Pe�᧔B�9��v�C�2<�f�GpY_
ӆ��͙ec�+	�h�o�<������xQeɢ1� OiGtU�[٬�L��i��k��F���/S2�Ϸ -1�����2��g�x�\��6 �*YX�ni�bq�:�����&�o���Rzީ�|�gH��~"��m�R��?O­��,-*4��P �H����a3Ͼe�}�������	'X�:l����kpu��S�q�g�m<���q�Qan�VY�����s*dzs6����{ �i=9�	�d�Xo��UIC�+a��{;��d���L���\�"��Q��,���fO���Y�&!��aD*����m!������,Dx�dp^��c�����ng��Ew9�P�x캮mx:7��c,5=+����).�ʤ٭��i�/�t�自�U~)2+�_�E��PVF,�՝�QC�m�����Y~4s�f,�EHY��]��=����T����z9z5��4�����F�⣁}�:��a�>i�t��DC�Ǆ���R�z2ve����9jqg��������Z%6j����?D.�zt��C�����s�kuOS�jmP��5P*: s
�,Qɡ�Y��<z�����׿чt���ڃ>g��6��1-#p��i��4g`������wBRqR{�vT����y�m��'��
rJM�W�Ɍ����&3�*h��y;o�Q�OO,U��"D7H�/�F�P��T��":�Ǧj�
+�R9r�?���8�\U�.Lf ��2\��j�Y@�n1a�W��^jq� �ht|~̈́ݴ�� /�_��,�fp��%q�ԣI}�_|��t#���G���H�6no���Г��%1|����RxP�Ȝn	F&ȒyL�x�hV��{���2<7.GG���̨K��ni1��b"�V^C�	�g�9o�v�;/�\��>�������V_�{��q�?1�Z0����������Q���ߧ`�A8���\g�z!�!?P�̢pÔ��D� o�hX�:��q��m޽c�'�N=�b��%a�������a1΁��:��/���2��a]kL�*��V�ݣ�.`2��H��V hz�b��6j�C���̐�&eE���)���O��a�Rw�6m~D�P�+vҢ�y�"�*7����r��Y����C��.�	_�������>����B����9�@:�Ù��w��K�ն�1W"�n�R30�AG���Xq�{%�X�e(j%O`����T�O�$��9ʊ�I��q�V�á�눮܊r���bdd�?�>漧��)~h���<ҁ�P�K���C���$Η���g3��g���%7ߜ�#�Zq��l����;��@~�A������
�R����r�NZD�$�Lϔ�<�;��Z�s�,LT���k�O-kib��4�b���M8���~#���d�OGVtv?�7΀�8�֊���A��-�b�3i΃8옋6Z�+��L��G��64���eŠwiEoY���j�8�f%#߸`�w���ަq�� �S������6p�6(��V/��C���?�^�B�7~5����$Q�m}�R�M��QV���0h�PF��"ZT��N)�ǃ r^3�|��>�3��\�����+[�-��#d<s[烚Ds�mJ�a�����
��d��ُ]7a8��.G�����%�A���gR�4�G�����S;/��n�+��1��kΖ�K��2џ=�)��ΰH1��b˱��hx�*A�dC'�����Z�x����ᢑBD�vVg:����j��Λ�V)tž^��E�HeM��;�![�����)�E�Hin3y�07O�L����ٲ^��q	9 ��{�u�YRwl�I`侘b
{o�zu��N��L��k�s3L�МpZ�&�� �3\]�9����m���p��H��R��re�)<J��0�,�)�pHF��D���c��DͰ'a�xM��^���_�Xr8
�Tf�����n�8e�=yQc� ��{�Α�%�r�nICm��sE����D�%�*{�!mV��Kx�F��	.ۥf����ite���t�d	K9ʍ�w�籡�Yu��l����	u��:#S�s�KB
���H���	�Q�Jt�h��X�CK��*.�Zb�`z{�/G^�{��c ��y�Ns]S^D����®O*�!�zk,����@�@1��0�POX���0V��R$�P������H���1���0B�2P������mnU8 -^���߈3�@پWM�T �+Dip����{k=�� �$o�0�$��P?��@ɚ�7���k��e8j�����1["��ex�a�â�|��Dk�N���y���p���:�#
���c����C�2j'=�wOۿ���|Z� r��m[�`FV�Mf+���C_�}n.Dg:�t���P)��4��|ݗ�Q3�u�,W^�N�>˥�4<�����慊�[�n�����M��?;j|�`T��vg�C��_�a�?$���lF�<�ɕD�1��o10�Ki6��.l@4r�}oJ"^�>�D�̤�c#�x~�N������){��o�#��a�iof�C���j:��	��?� bn��9�Owѡ2'e��,�d@��{:�j��dć�%�[��w�Q��Ӎ9��j��W(�e(�R�}wྋ<)�&T��/a�[�i�<����Kn+��&����չd��0w���B�U��6x�Q��>N�w\3�́��l�����w�����bDQ�{�7�
R`��ϡ����~��*���a�2"`�>��~���@~8��^];O�
�u!���mi�o�o��>	Yo��u�H��޸h�KF����w���N�r`Iן:�QGx�ޟ��D=�l�y<�\aE��Q��T樍�!����F�25k�U��3E=�p��?]?%�P@����R;f�K�6���w���\o��G��Q���-���.;F�뽏+0P4��L�o������Q���H�:���V�տs�lZ�ǫd�[si�%�X�A_P~˪�*d����̄`Qv/��A^#���b�b�k`�D�P��ݶn�苫�x#�q���	f�܂��J��j��z�L1�͇4F|��5�ǜ�h�ej��a�����u�@�5 �3
�g2^d���o�_aG'Ͳf2M�`գYN}�HY�	�_i���U�Z��\�-Ǜ�O7鸾�Dv���"����?�5���(:�=;�p������e.*�d����zj���D�p-������	��`a������nė�!�Ϝ�'Ѕ��$׬ֶvRxS�{�������po�C+UN?���1d���$�E Ke�t��@e �ӷ�EZ"H]��z�cc�����:wu�d'uy�at�1�/�s,��G:���o��H�e�:L`�ӕ��пx��w�m��7���4��h�s^�a_������k�\��O)��WU9o���2�#lS�Oj�LloJ�~����*� E_rbHsz���M�s����<֡R����N�4�M3i�S$�yM���0&�_�@d1��
��	%�(?�����>�e�eG9��B�쵿^�}
����Ĳ���m;ѵ����Y�k�ϓ@�|C/�=QE�=��J��	n��Bq����C����S�n�i�d���������^��e�+��9�4��3��D��Ʒ)�1��<��[�7`mD*���k�7�bz�J��?��No�͈��a^W��eg0��b�j-"����Z��W�A�Q�/jQ�2
N��I.���ӳ�Zy�]���1�4���ry�/q$I�
��8\j�~��ŹkN$޽�F>?Z���%;�ځ��h�V�u�j<ǌ�Ib^�q����AV������ŝ�h(�[�u�Rm�PUrA�)`���l���pxAȳ��Α�̄�@N�m�8O4��<�����ć<.��c����$�WQ6!+��
�x/wB�.?���}m+F��ݻ���|�����RwjyS���_K-R}���^�b/Wm�1:�i��/�p휙HӕA��qO�wh�Y��s�@���'/H7����%S�\�r#���<~J�N��X��9ShV1�,�q�<�$���XB`w�5Z,[:��ՒcJ��eD�*c���ά��-Td/��=�^�)����Z�^x���g����Ii@�ּFa(?�b8!��a�R�U"�]C2/��?�� _N���{柏cIa�����gP%�5�	:ZS��ׅ�'l�f'�q���D�\��~����o����Ycd��ˊ�w�-z������F���>_6��?����\A�̀�y¬ho|����$�i�>2]ؐb��]��o�� �/�$a~'�'���XǤ�F�<<�/�]�x�Ǵ�_WIh$�����筒8��j.�Sf� �pXW,���@\����1�M#=V�>��$Clu(~'j'ũ��@�s>-e'��z�i��}%�vRA�d|05ނ�'R�M'v/��4h��� c`��x����~(Êp$�]�W@,X����!�t��[.�މG���9����m?��T׶Ⱥ��h���jp�3W^9,�Y.*�i��=1qP&.0�I>�A1oR��
ǝ���+��t���% �7����	��B>U�u�]l�?�h�P��ߙۅ�X{�ڤQ��Q��tD��m������))�k�1�2��]yU��[���#���c��k�:g�@,������f�稊S**����FEA|�����V��b�!�,kV�J�}��Y�(8���A�G�������P'�&����J��6�°ꝋ���K���c�X~0a�eevfl�o(� ј�=|s��'G/���N�j���g3 �-xu�1њ
�y�\����O�G��@J|�v� �Cj>1 VN1[%w�f$m��������%2;͙�o�z�q��ZS�[O�D��?���������Q��-2����bPYME�W���ˮ��χu�'O�uΧ��r,������ͩ��.�ޣ�ʑ"e���|�~IV��$�U��%�6���t
���8"_;R������*x��Y��xKe�º�35�X��ܗ��h��� !���b�ZU�K�Q�
/T`���V�ISVG$<x F��9_�9�N��Qʀ�3�]�����9�7}/�ɷ������6)^�J��43d|Ԍ�X�G��	������#O۩����{m4��/�����7#�g�%Tr���i�$��:*|�4���fI����c���R�㟗�i���,�w���{O!����B�a��~YR��c֥���MC�U�b=OO�噀@�I����	�*<(�t�C��
0�R��N�(c��@'X W
a��	C M �_��A$U��vA.�8�s�b�|Q��X��Ob\VTE�gqן�\���\��H�q�gjQ��V�cʹE���6����Wo����PAh��;�t��ߙۑ����cp���C#���z,)蓕`�a���͐^��lO`�_��Q��i��>LMyo�]��gR�o���*t�K�
�x>e��ŏ�-�~H��o��9�3Fb
��Ճ���/�7�tB�	c����)-Mg�}��K��j�(��N�n"U�ew�C%/|����hj��N�嘆r�����Pa��g�!��	�H�E̞�%f�� 
!� ��{��Mo\���Ѯ��N��0{Mz�����t�#(��+��K�c�\�K����+9pU)9$/��uz�0+�����p1b+�!�#�5����EΒt���o�U?��f=W�i�S�[�Eݣ��K.��2��-��}�⓰>�z:!}I�m\�$�Mpzfpg� ��CXn����ߵs�Q���m���������sf.J �eHPS���Gj�C
���s�l,"�^�[i�63��.Ո] A���n�S�Z�^�Y���u.�����C����B��o\uI���"��@OQ�q��1E��|V�b^�&��S+�Ͷ�����L'���n��^���$��h��)D`�~N\��ˏ���)���U��ŇZw?��{�����L��E�B餢>d�}���9*�_�g�\�M��+��������S���}}�ST�LB����chG�BycT�Ą⾦��u�V?,���^"x�
Pm�A��1z�&� p�-V��Ǝ$�_��%�S�s����:@m�8���.�['*͖+.��v����x�W=�d�+�\������V;_]�Kې���̠�=�OZ�(3�Ӱ��9��3�R'�̈́?��O�4pix\�|�=Β�$��j�9L�Q{z8���XkR��{�j���V �=�5���F��	f��'��K��P���念bր��@�L��؁��
3p��!��.�9��P�·/䆖F��5��t-�9`�;��\�E��_)��	>�.
/s ���5Zt��8�l��$^�0`Xy��J+`j�*�4���ߐO�h��J���PY�d��)�5��)��k�zY�Ճ
 ����iJ�{	�*P�2a��5�pʢ�"�J'�6<��LZ�� w���!���r�ݰ}�.�\j>�bZ��A[܋�C�.ܺ�'�Zό��Y���hP�>֜��f	w��jy�]���s���Dso흔n�?�/���&����D��[�/���b�-����L�wӞh�VPx�-Z�׺��0��������YN j!3� xw���r-�Ǽ� ����0ENc=��(��[ ���D`u��u����VU��p37陼g<�ɕ�HT�M�Ij(-��n����1�_j�GeL��v�Nc�f�o��O;{�N]�X�����_& զ�.w�p�����)�Cc�+�v��Y>�P>/oX4YDlt�Cn�A�lP�����|�Z,��x�i��ì��t�bqe�ջn]G���T�*�F6�fr�pŧ��㱥�g�����v�7�<��y��sj��l�z`«-x�s�*�r�y@!���2q�'J���Rl���5Qy�̱x���-%Mr�|�}g���_$ųN��|fǗ��Ri�N���V�
j[��'v�����h<����ߤF/4�C|�7���4��mƌ��6&m�oڽI��y����xW-��7h���q�]�o��Ƞz	�@��aJ�����X��ù��+���]fe�[t���"�����O7[�Ա�>��q,5]*,S.�<���ⵗ��
d��1�?6\���D���m��S��B�9�9O�-�Z�H�o���AX�7X���`�K�n69������\Q.+Ga'��sgd�xk��QX���A�a���"KQ���P����5�bp�
)U�"�l�7+�da��
,�\���eO�aQꏑٸ]f�԰��̀�kv��k�\�TۅnL>$�4w��<�ڐ��� �85��$�Kb�/�s���bR���~��Ȯ@e����fAYVj��f`��4�<�3�90TS��.ߤ(`at��^Cw�=���'+I%�x\�xgs˞VWm&���¾h�j@2��������6,�ǎ!�8o	����/,潨zظ[��sU�W�VdҼ�aB}�~� y�\O�F!L~�x�%r 8�y��.�d7��{�v��;�3n�HD��@�s�����n�
~� �cV���/e��eѠ��
��?练�I]Λ�8�rY`�ڡd;�|B��Ы�X�*�p".|1fZ�[�y���?%�3���-(�t�M[���yP�\@� �^e�ީ��@�*8���a���O}�z
��@����fOM=v`�O�˛�`��5B1��JhY()]���*�ػs��MK͉�4��#D$:X_&T@��7�F>{�kg6.)��ua2xj������EG���R����������>{��>��D�rÅ���Z)�Ug�ľ�K�2��G�Ԉ%HR�O6�\�;�o�o�~\�p����#�t��������?�H��=_�Z�@&B�ʇ::�L4iO���^�Vٿ�<7kZ�o��U*�
�Y�(�D�.Sh91�DZQ�'F?�W,Q��^���-W��[j~E�'0?�%�p��`a�Y2��%e���y��;!(.�nY���4D�XtcK,3��Ua���~�C�����c?�D3H�ڹ4n����l)�]��!WQɄ�f�����ub]Ge��<�:Q��e j�y!��@�R�����b����y��B[�d��O6�J��B��p�uy�-ة�m�^G{rrH�a��~ןm)�<�טu��-ÀmUO�����'J�u���ǲ��gçi�F"����9*����"�L�)���ɮ�(�yζ��R&0-�i�)���>^����B-<Mf]_�,8�z(/]s������1�X��]|w��w*���6�L��
;��4�J�y�]\M�{�6a=�J�����(��D2l��W孍i�?�d˚�MlCU�t.b#
�{}� H`D���9���<�ge��-\�iL��CL�r��b���$����WĹ�Yj��_F@�a.�h%3����^����5s��q�����/I�Vy�\&�P9���>�0��e{ᬵ���[�n<s>_�+L�)t�'i$~ i���ZI�)�z�:���FzC�ц�NY�r����U�+&�\��I0��Z�8r�\1(��,da�+Y���zF�}8�y��n�
Mz�Џ�j*s����$lMiQT#�=.񿣁��6�nW��B����cډ����hPZ�����1����њ��rw$�Y�*������b+oʇ�d��Lը3�ٔ��N�F�"�Ux��.�%���-����dҩ��@�c��pD��.sJK����	�M kz#�;l)�+;A	����ۋs�7�(�J޽a��Mvb�����6�� �ȸ�K20d�2��nT���E�x�R��}��X�5���P�v��U�M��(0��mT�!\8o~��H�D�<^���eo�ЌQ�6���,E��q��sg4���Na�� ��D	���ѥ �ѵ9Q�R=\4��nAm�{�3��$lA(W닣TS�D)K���E' _rT�%��r�?�m�&r\Y��n������܍�������!l9�_�7Hj��~R�&���K��Q���@�KH��D�2[�Z�	Fl���E�U�,vP��;�������^��PW�ħt�g�M�}z�s3�ڥ��vu��a��(�vSx�=�Ω�#�����I���4�!�OA��KQ5춭5�,��
J�B,�n�W�+#d�K᪙���Z�ߘ����G�-��{uM����B�Ra�ntۈ�7|V�����Vۃ3#t�kk�����-O� $2��#�ę�I��[���ǀ7�K"_7��4��Q�e����N ��	��NTF�BA}j�+�
qn�H�����sU���9�t؄j�@��qeW�,�	a)�cx�Z���>��Is�) �v��'jk/�q��/�7/%��ۂw~����:-��{�Vc�ҰZg%)��-�m����>|x�t{q5��|������Mӏ&���샂����Y� �צ̢ @�-����w�| ���.��]z�G`�����p���/���/d�b�z���
J��g��Ȳ��]įN�y6�����2D�G��Tvp�H���KQ�����o L�
ܢ+�h�ˎ���������� ����V�/�Y�svP?�J34�|�P$Ly�{��uJ[���G�d����YC���z�Exx���y�\(�%p�n[��l��*��SP��]�1J(��R���fu<�^s��}�]#&\������Q�XI����@����@�����RF�zdy � x�k'vI>,F�&5^��m��0`Z��>9�{��7Ne��H��c�"�ݪ��nZ������{�V��߀c?&v2�_���Yq�����S�\Ɉ��C���q�B���Vr�P���¸���AeT�g�%H�q��|��9أ���u�D1H��4
�%H�S
�д�w>Zpl[���.�'�ֻ��Y>���+���=���>D."�2�,hǃ|M�6Ć��\�,'�=N�s�A�о�,r ��,,�9��O�4L[��?^H�~(E�Pnf2S��g����i����I��R����t��k���cm����q�_���X�u�7������r���b��.���G�f���\D��+��*s�������Cϼ�����jGQ@�`Ϣ1�<��i=Z�;���.7��c��L`�<�S��!�KLpP(�n�c���L[�b7K۾#{&Ƈ1C��IkX'�}U���<�Rke�a���ס����9��Ol�����yTI����8c]�\�BK3{F͹X��||m�0h*���TH5s��[���"�[�a���-�%��r>'���-R�&%���71��k�I�T���R����5���:7���4d��"cV�S +��e�j����!���&`�ǌ8���у
$�p�oض�k�k�1lj8�m@���äy\"�Y�S������s#�b=-&��P��[�*�|���L���s��y�A��G�2��ݤe�?�zR�"���Z��䭞���H�2��)Y%��.�F���Y)@R�9]�op-��E[E����K'���u�'��~��i��b8Ξ��XkB�J�`cFNNQeB'&B���QUn2�����P��� SCim_�@�s4R��ϗ�G3�?�@8�)4�%�n� Ċ�L
�@���y��_�;���7�BL�g�Fa��L��>��rK��L}s���v�s")8�zf�;ѻ�N�n�ݴA���\#���b��7$ �
����\����~4r����1��f6�0�ca+]}���ߗ �y��ԃ�O��C)��.�Q�6�XHz��l��RB�)P�E� `/e(��xy���k�r�]�({$�M*�V4��th����-�Y�[��:@��HDn���W>���r�]֜�<�D�[�/��PҨ$Am)����,�����ϲ�>Ѭ{n��"+�.@(��p�C�ȋ��V��䮌E���*��ұ.�&`��w����
g����&�F_���ӝ��E�6�N�-����������6��OH�+W��&}\�u�{/r�u1U�]�C`�Q0��k<�W���0�A�YV�;��s~�-G����j���TY��H�z�v9-��S�C�=r���SW��Ӥ,��̜ݯ.X��!:H��9�����ۚw��ťG^�kG�|���5�	R�����Q�$ӏ>V��oD!�n)18a$�m����a��x������� ��BA�|�Ië��_�~J%� _C״���G�ȺW�n�k���4���J1�4L�4�(M��K"�B����n�1�L`��T)��<�o�l�Z�h�#�8 @���{����[@�{���uے��J��FЇ|�o��R�.�ҥ�M3F��m��&������|~�	�����fys��O�g%Ҷ����(Mdd$L��E�vP+���|��QՖ���K��6�!�_9��'9�]�9�~5��VW�{ ��.��kN6'$6�Ę�����
�����m�PK�FZ&�­]˕�6#�'s���q�%t��A�p�%���:�^������!=#ʎ[H⮳�C,�-wB޻�Mjo���:[~�Y4}T�~�3n{ ƚ5�!��5�}�_D�����C����H�/,6a��$W����i7SH�n(����֊E;�Ԉ�qX&��L��"6*:n��8���
�z�J���xH��e�������E$��/�H���i;X�0U��wO��ĸ�$a3"�U͓�� ��3R�l�v`�q;?.�i͝���2iR�I�$')?L�@�_���G�z������aa7�C�À+x+2R���Hg؂�|��:�i����8��^���*/"3��#���B�Z�"KĘ�?ƊU۷-"��M��������X����f���*ϩ�������K�����0���^w��ayH,=$�f�ԡ�
>�5:Xx\%���t���Qz[�;�N*�Rai8o&���iL�����D�d�b�U�`<���:�S�ޱ�����Țʡg8��4��2�!��V�ǡH��^OB�ML�R绂�5�]u��]������ت\�t�%&w^m�e��
Ç�<1�Y�F)���h�׫��}y���=f(v�>�44�E8��0d��t�(�����^Q�V�o������b�5��H�[�E�oBNHA�%˺���|��[>��[C�w���R,�B.}e�!7�d`�ճs���G7X�=���s���x� l����qƘ�[��H�rS�TJB,<�Ō �@ ��ݻ�9̝vV���[c5�CaR!5���t�a��<Vi�
A�=���e�� �
���U���})�S��Dj�b�@{�$Uw@��j�g{�e���U�/�~Z�^�J.B��YY��4Qu-P�&��]�V	�ҍ����q�ŏ�~\կi��xVwIb>���8��s�@&�ΆnX�8Y0j�������nՅ�n|�5�S 㝃�����=���D0!����lFm�i�Cr�1_.�SE"������E�ّ�
�gH���d�I�@��܌��}(=SUS�܎�ͨ���o&+��F��sw��ӋR�SF���`+��rrn��;�YK��Ae-u��1�+�m��L�-�Sָ�5��)����<�X*Dd�I\D��g�~�<����s�<��U�;��E��J+����M�NY)�C��G������ċxǡ:y//���`�������X}�A�6�Trb��|Na�$�6���"��,xZ�5-���>�pmM1�C�<W��T��g;�@i^GR���6���T�>��x�I�%��c0l�{�7����6�4�v�9�Mo�`��.c��.8��~������)�L��|�}� �zo뚫=�sBw��
�[U&�v��,
ޅ���q���Ղ�-�އVJ�Xxe�d�k��͕��$n��+%h���㌋=����XP�~>̰���Y.�����<�,��;fEN�K����k��J���;?�$*Gо�3�+�_�hφl�!�l��2z�
��Ck�I1�%^��6`럪9;!c��-
��LU��Y�j]�s�~�o��Vn�Ah�MO�7�_é���u8m����<��xQ+��X��䙋�΋��%������Gf�E�c{
O�V�[a ���j�L7�$?h�骶k�`��(>�\�Z]�����3�p�k#A'�ҍ}�㨞�����S�����J�<��5\�(	ݘ`����`p"h�W!���g�:'�����5�4����875�t�J�!X����5lUL_X!+�p��s���6�r�S��]�3�l�>3���a8���E�ɫ��n�Oi���a�9,֝��(<{	�S�ч�=��#��<��.�k.&���&�(�������{ ��4�턾�n_����I?�Uy��b���u]Yp�qk�N�&Vw��#�o��~�H�&)P��<��kA���=�c��4�B����=D�@Ѐ��Z
�>/Xt6�ԓn��0��ס�2V�Im���6Y��zU������S&x�g���� ��x�j�ck�/
�'���B3��Q��er$gYzM�� ��v�v;�-vҝf�0���HãO�
���kR�E-������^g�9c�s��S�nO���a���D$"��ܵ�i�!h�
�Ђ�h�7����ޮ]Zj�p�|�D�z9
��*��L�G�2E�(�A��t��
�A���f�0nF�g���28ͪ����L|�)]E�|:����L9*1����Q�З$!l$�ːAr"C ���0������{x�~�m����R�{#������<�F�c��u�l�K}��^"��U�y���Ug\��w�'���GQ�e�f#���7X뤲D�۴IMu�����q�:���˺��n	�7ˤ[�Ψ�&;���J��db��6V�����&y��F<�
�8���綠�m{�`�Y/��AL�'sC��t�`��&7�	1��߈�1"z�W��V=��gWH�N@��<���Uϟu�*��<,��t�#�����n7�t>�� V艕t+(2��s-o�O�"�o�p'����7�1�;K*�l�Йg'0���餃v�8�0�GH��Gؓ�$,)W�����d����u�[!���)��Э��U��N��+�/��:E!�Vv�Fi��e8�N˺�-�b�Z�#B �D��ђ�9���²A�,: �y]�1�s��"�(��U��؅ӷ�nW�?�e^jYO�"�.��HgO��~�ت�	�\�|��f�>n�ծ��Jس�`�(/��@^���z%_���b�
e�q7���Ĝ�w�/����m�����3E)��UБB�_]���6�$�ՏW�%�2������]ϖ�?�P�	I[�v��PE�[���d��1\�KP��шx�澗|ƭ��-�� x�`;���zJk\��6�����b�	�Ր�$<�XMI�͒!��?�|��3ON�"��nò�l�f��~	&)�6.~�����<�e��pi�;2���I{���(��]��A�L0���S�$��!荸����7<&�G��iF�� z�~�Ԫ���~B�P��k���۟r�-��x���!����^��,#rJ�-�}iG�XS(}�\+ �;�v�����L�Ur��7Uv��r�
���aϵ�4 qYS�C�b�$Ο��U���3��3s	t��ډ����2�υmO�\b)J��f?���7��W���*i���eu$ߚ�w�0��p�&����`O̬(���q<N@�r��-����a�5̯˯�Շ���x��^�/W׻ҏ�0_m�+&�=��w�ltH���z�b���J�#CY^��#Ք3�&�V4�3[ۗ�շ3b������e8�-U#ެ�^��z��
_��[��-BP[�x"�ƶ�F�I�*����Qqj#��@؉zP�| o(=(v8|����Asz�a)�ݠ�G&c��\�,Gq�������H��v��G~��J�Q��XHd��)̎�|��o���jv�_�ixq�����8��G�p��f4�*�Il�{J	�8c��9eH�\����ԧ�ߔ�m�O9��by���ռ[N�f��a#���h[^P�[�F�W2� ����8uҘ�Z+QR3�r�3��������p�]E�UzX��4���{�� R���V$�$��H�t���wh"5.	m����V5֧���N��\U���d*^/b�����5��ȳy�G�-&o������%%/������8��H�U�,*����n�(۰�y>d�&5֒vr�ΙOh3��P9���oe��Ri"!���a���a2ޣ0���y�EL��Wˀ�G�(@;)���&4�`��"�p��ё��.�5N�&"�*	O��yA)^�q�tч􄌁��i�k�<��0U�-YE
�7���*a+4��X�C����P�,A�����'�E���G��V������qn��Y �T.-4�t���J�d@�w���%4�O����s��e�w�?���6�77 ��E1]^趉tF����0��N	v���=Xq'�X蜬�3���J�o���F��O�A���g�9a�������NE����D~� RcMWi'�|�p$A�����&T�R�y)x/e]�����O@���_V��#z$�Ƒ����\�3#���x~�z����7l1�~�\X=�|o�nQ��@�6�S�dE,F��Z����1#�t��`g��D������Q��}��n�Dd2Jzh��������Ĭ����*-7����_�6���h��-x�i`�aχ�0��WH1��W�sX�3����������̴��v��c��]ݪ7Z��`X���pU�a�i��X�n�q݁��	�j��t��� �;�bsҁf��v˗RG��/yB�4�,¶~��  ^�l����%ov��ol���������iF�����9��@�#����T����D���g�#,��'m}ƫlS�&�S�X�2޾l	���v(���0l��j|�4OJ����3ϲ��F���WJ��Ԝp�����[��N����9M��X\�_a�UVA�B4Q�ȭ�H��x�R�ܓ"�R����&����U, /��U��5o%��+�mx@�����&��}?	a!@[�OL��t�^��Y�P4�]P�;����}��u���2�(;��0/e^(�i�m4��������*��D�x���}|>Ө츰3���v�mC��㥤O�� ��!a'��EM}�~ŷ�ZԤ�d���J�)�� 8��x�`H�����'s����i��=8�
���0z���l)�g-���#p!���=^3�X��P�#J=����
�|�F�+'2�#�F�n�m|R�2Ö-0/j��n�r[�����+ʾZ&��8����E�3f̑MCX8�8�Js\����x/�Q�ø����5��K՟<Dv@�ˬ/�!�j��<�B�9��nX!aX��jE4��
�Y3�F�gWJ�}�18��`�(LR�QK
m��T�m�YX�<LN�*�[�0g�!�D�Xu�Q���u�#a<5���m��%#_ŗީ�[m�.-�G|�����l#����������o5�R��	⿁S���!�[����G��X��Λ'ߘv�ܖ��#W���6^�?~�p&���-�Cĕy�)��a
��)��aw�����\���Q�*��(������qG� /���%ϭ�]� ����)������i���M�0Dp���ETk^�3-��M�bȆ?x�3�;�"D�J;�y���d<�>Ħk� ��7��YK�M�q��q�����������nQ J�󬥜̨�� �oZ?L�53(>��=�M�-Z@�#�w�3eY5c	�Q�?m-���5��Q��4���x���|)@l���	�EtI�n�d(6���Hy(U�v��܀���G�	!fez �1�!�=��٭��!� %-O���K�i�e�@궕��@�d"R���C
&�\�q��((��˂�?�N���'�w>ܵ5�O�����d:l����kZ�:怷��r)��/��,4_�m(�8 ZD��>&�=T���"�u��WT~!�d�qP�cp��.��ZF
w��{�慵�����o��#��M{}�,M�2���]��4��i�WOL���	�+3�taɷKR��d�<��?�8d�^���p�z9fhGC	.�*]8���Z�_��R!zZ
��i[x�օ\��F�.�[�1tS= �����w���F��Zk[�����X�|(�X�;����[]�L�DP�Ɛϰngɽ9;�!���M��K���Oa�q�6��TT��9枾�J�/::
H�֘P��^�W3t�� �=�3U�ri���7�Uv�_���lT)�T}.�J���U��{;C�D��Uv���a���W�#��"�߁�w�.�>FpI1�h|�ꚏ5Y��˷��2R��QB�	�c�����M�NȠt�E��J��{y�".�EU=n��1��� VT�j�XD@����}���Z:A`hmH��"`�M��e��.�`lH�3k��;+9A(0��X!���1��o��m�:DvU�s�cY��S�!���hI�1	Q�N�uQO�����
�;��[�!�ٝ1zFQ���o�3��q.�4J;@e�v�+�g��	�sM��A/�����<���G3] �\�L�9�)	s���?Y�,a᷀xS���`]�t#������ù���(va��.� ��
�3%a�}2�N�� xTaX�0'Ǩa(+@��q!��S~Gg���`Q]��Td}Ic$�Y�j��anI�sQԠ�Ji��z��Cs`J�B����SDp�pK�v!	�"o����d�Z���$�6@k����Ԗ��l���K�Δ��m�l�U�F�m�[=j�Gm���ix�g(P%ͧ �Z<��{a�	t5���O�k;U��qٰ�h�$4ۣ?צ��u��[�R��%5�@c�5H�6�X8$C�ă�ߨ骘v!���i�H��fC��������y����_l�w���<B"�W�p�B�O���4��ra��]@o� VvIr�Tw�5_6[ߩt�fI�g���
e2G�{�d���?�_No4Q��"l�ݨ�7Ĳ���}�b�M\H�� D��Y �'3�IwXX�|R�ÍJP4ɷN��PS�1��2���ŽT� "�M�*������ �K�,��G��`��}����@�2J@�#�S�x��;��N�@�t�T��S�[ra�u���xjם�� �_�+/�*=�ᑛ�kL�[l*I���p����|ׄ��S^�Ё�l��6�*օ�c�oF4氤d��>���QU����  �^[��C��/M����1��D� �'y��?rJ�$~�9��^�x�|1�3��A���!!4�/�7��B��Yqŵ���D�I�M���0��7u��<x�@��R@u�L�L��䧲�!(�m?���e�{F�a������x�]V�y��2�s�e�!F��5 �B(<��mP?��� ��w<L4V~�y<��sѶ"�G�i��Zr��N�CÈ:��.~�DM�`�^�<�~s�����bV�I".Fn��ޔ0�0��V�,��49���b_,`A�]wI7�za�=7�!�B���ll���������)��'�?3@}�$��>���I�\�C^��&���ӘApϨ�QKH��F �t�(���|�q��kVJ^�����9���U�1Tp�rP����j7��8���LD\�h�����٪��j��@���p��k�ve�Q���&哣>�r�;c=��8�'v�,%|����9�	��?M��y���9���yt���I�I"�|H�ϩy�$T��/��~&_v�M��{	�[�(�M�cц����%I�ܴ������>j�b�g�L}��*�x�da/X�a�ʖ�d�]���5#�4^`h���p"B��D��I���4�c(�A���h�m�)�ԦO�I�GITfr�yR�7օ���K.����E�i�ψ!C�3�VE�X�o��|aH	W��Hs=ܭ�NR80f�e�QUz<��R]/�m���Å9�4���`(�9�a���O�&���p��Ħ��`�5�F�~�j]��I_�V�������Mig���T�r3����R�UR�*p1������nN��g�|�}a!���ٛ��afot0�}����{�h���"�ſ�b���ަi�5�n�`0�p�2�d?u�.���=K��re?_J Wa�<�LO��ÂY�@��0�?#�h����$�(;u�OT��� �c�}��惸2���N�C��^�0�D����*�;� oR��IG�Z��!�/f����m����[���l��uV	� gJ�FEN��U-��&��A�z�]R���\�hii9���G���̇��|��B��yw���U�x!h`ވ	�3�ׅ�'�Tx^��vj��'j��,^�t1�p,��zc���ʖ�_x+��@���d�}5M�%
�z���Ο��,],k�
��W#+2����g��I��---���L��� � JЩͭ)�N�1�`�M�؎
#,HXBu\���I{��
:
G"��l�2�N�X(�˪� @l
s�.PY^CL��0H��p�yd��K�)�r�e{/5w��o��\*g���mI>{x�gٺ� �<���g��X�ۭ�d1kP������9�u⬅����+�������?��9����a�0^vώ��	�k����Y F����K>�f��-m%Ŕ�����ɗŝ��'<��󱾢�C�0��յq+��y��7�"N�b�O����N?�sDFG�*�@v��}L�����m���u�d�W�ta��2^p�p8N�J%�FN����J{�RT9Ԥ�cؘ��N�k2�[
��6����Y�T�g�1$�*)�����T�����\q���ݩ����p����Tr��������þ��&KŹ�����6��L�M���*��|{��W���\Њ�-���^�YV�tÏ;'�6ڿ@�8����3,�}��#Ϋg9�m9�$�G���QɞP�Dd'\���=��sb/��4�8���A~z���Ba�+ةu9||A;9�  qݽ��Z}��x�蒀+ ���Ve%�Y7u�z `sx�'�6��K�W���t�-�o��$��Û�^� !�\b��`u���p�Ɛ�Y
�43ô�<��k�+�a�ms��-V��'~I�OX�ӫ�5�4S���ViIl.S]\��S�K��꼚ST����*�y��cE�I~T�tE���OW�%u4!�e��9��⊆P�\���{���#�}�NG���}S0�?�ǧ출��"��`K�k��6���:�uS��6�X	�RR�I�B���6XM��6[o:����C�4�����OP�rZ��� �8=� �ʦV�
�X+X\,TS-0<�
?d� ���MV��d��7٧�Y&q��ޠI�Uqk�����
�=i{D7Q��\��{R1�H#������Or��sB�s�����ɭ��tr<)~����%Kw/:�,�d
��G�]���.>O����П��Y�^���KH�ɮ4�?�&���jSԿFz3�E��ɇ-�F[O��g��we!��Td�>=�u+��n��H��4�C ��{m}�̇p�LS�kk�l}��`�}�'�=��v��z�$��c�?T#����]����ϡ2���;�7�,b�DA����'��(�N�B��#���-=V��U�0u��RR� m���͹&L{ 엽'"F˼{C�#���/|�ފ���ئ�e�4�� �I䗩Hq+]�����x� �_����!���T�}$)�+k`�e���
=��^��Y��
����4��?�	����C��x`�m�ޱ��c���	.�oe����� Yd<�qgK&����A�s������-n-~�$W�Ϻỳε}�W xw�1�Ne�k`]�i,�;!�Z��Jw�?2g-��h�����ů��dch��Ѭ��Љ���$�O�tXк?�6���N.J������c6ED�DI���cN�� <<O�e#.��]O������V�7�����_h���?-����Wb�h�yx�~e}g����_�[�)��*uM�0YW�&�X(���+4ר#5z+�Lu���@�E7��Xs���S]I �����{N,�k�R��i,.�+$��X�:�8�� ���1SU1�yR������`�Z��Cؑ�Z*�Vc�F�[-3V�n`.�}! ���DJ��Ž�xۤUeE��~9a6~M_G
�.�0
���� Ͼ"�va�y'v���,���y��6��b^�6P�M���3=#��jWn��fy�0�P���QAsAܠ����ʾ+�ϵ�5�d/���r� �#�,N ʖ~p���y�Џ7TS��빯D˿&Hϗ��'=��h��m��3��M��~�!�*3��V��צ��z�6�%J������bu�/vr:�S�nj��Z���,c)ӆ7c�j-�����ݥ���Y�bV#>�r�(u��&m`�[�\�	����~A�a�?�2�=�=�J1s�d�ͧ�P�#z�u�p`t�w��]��+�z�?��أ�
��W���۞��� ��4�5[�Ț�(�iW���3��$2�9�m̢��݋�@�K�~%3B&�!�i�S[`P�5�ځ4[p����z���Ք��F��H[�=�c$$m�/��+�TH`�*W�b����k�[�T�k�[���䮎�۸��~����oW����)��
�"��ƴ��,B��l����N{-�K�q�9<ߥ����:�>+�o���>��[���T�Έ^U<�4O��ˀ�\u�g)ź�Ye+ �94�#v�+S$���^{�l@%��:���e/�II�Zq5�D}��G=a�i,�Se��oCN}�WH�J��W�(�y���r���,����<>�}/�k�c^ԫ;�Ba�d�m�5��4�b�a��X�o�դ�ir�W�B����S��~˒���v"7D���A�G���QB�iBrCՆ�&��d�X'v�VC5��jv�5c�l!��E�ͼ��"�)��[�^-��P���^=��݅6��!�I�j�v�K�}��򁘠�@5#�/|}Q
��+r�]®^���q4�[�'e�h�C���[��O�#�]sh��癒C��~R���R�P(�3���3�LiTc�{9��ꈎ>w��0��Ht��20�Iwٰ�(c�))��1#��=�&j5|��q�/v4%(�\h��q�߄�qe6.���Rzu��*1?}.G8v�Dʠx;J���)ɬ�5��N��E�>j��5��W+�~��и��e�o�rO�\�r,�Y����ʒh��B��p�#��ե꼎��EK*���݆�-�K2����@[ �dwe�CtҠF}ӕ2����_����{�V`���IRFʘ�rc���6_4�AD�u"΋0��8E�d��HY�pf>�NV�>���~�Su'�O?���Yh�{1Sג6�gO�,�uN��]P�}2>9j��1=�њp!)Uv���`I?��Q;�x�u*�.F�2 ����Bt�W�������#�K����in��HG�ۣd�З��a�5��¿4��/Pj�~-eU%��X������i[�&b�)RWK"a��>*���,����z鶱�=Аa�&	F)�p�s}��R���@ŒSr�5���Sp��tr�@5�� @�+�Jv�Nn�Ł7VZ*W�P�Tplr�D��G�X�(,���=�B�/ȕ3��@\��Y�M�����~�h���Z��L�r,�,�4bt����w�����N~,[�v�b�{�s��TrK��O��#�K���jp�a��:^�Bhߩ��>�G�Ik4�!/t�п�_`9�w����
:*Ѝ��)�!��_Ww)@@Ͷo�*�n�oI�![:���i���|��*q~=/�G��T��+�vpE��F�|+[�:c����
;���Y�ꠕgo�U����ػtQ��C��9�����<���0��T����{]��.�a�D?q�nEX�>�c$K��|FCI��j�NIoC욈���B�Q�����$)� &���ß��'.ʮ�ο���>�`eڭԱ�]��J�YB��Ôc�p����[��>�}
�~Sd�;?F������z^�)d�JRW�.X,0�Q�>^���B��6��.��Rlz*�����-)G������T�e���;����w�_�x`�C�x��f�{��!O���6�%�LW�����_f�>D+�Ӓ
�&�m���q_�G�0��R�I�2�8a�Mm��Ty<��}�e5��K>t�����
b�;PqMD'���LP�cV%Epaq9����)Osѯ��q�q )���O�%-�͐/%���$��E� ����[��I�{�ڬ��|e/ޛ�_i��2�[y�w�u�9���?ii��v�B_!����K�!��&ܝ��8�$�#$]��i{��x�/8���u}c&��K�P���ܳf��``�n�'tj��VT�I4ެD|+XR�A0��&j����T�Ts����m�|��R���������13�M�!.�/�R �*ŃL����tyf���VO�+�-�ח������͌B��T��Ns馏��1n�^�!|D�+eD�H��}m��7�P��hR�)((�;\��H���:�4&Md����R�B�#г��֔�Q"pQ�ϻ.�b��L�����mD�	x1~\�9�Ye��@�OJ����{��'�������o��d��ֳ�Z���䊢�n�]�z���o�e�0AC��k9�Q?lmN���\�_e�������O�QV��WS�sdC����i܇��`��V%Z���da�i����#H:"�;T���$�#Q��>���Yv˒�Y�!��� ;��[UT�AY�[�%-���O����]H�����&��=Pt�fdJ��=���g��[!��#���Z��:��jW':(vQj��B�z�@}�T�)�q�V��r�2���[F�0.�k�5'R�aR\�1���m�N���J�e��^�����-a>TT`_�c4��2�K������ߧ�sMO텲d�6�嬏�NY7�0p�lq�x%�72�\ϑR֪�%��D��!���P:m%(ڑ��B.AA!��7]-$m�Ԩ�H|�G�m~
2���=��w_D6D^�P�;5u~b��s��

L�IB�*+��Қ<K��;��?��{5�`K)�G|b�%W�-���p��RF1N/�� ��u1���Kf�;Ԏj�3�d��5��|�]
�C*��5r�/�M*���&cNʧUYbK�S=g��N%I���co�ʮ`g�T�DE�x��-rFQ�t���r9�h>zzanV��1�����Z$h��a��f(�H�eё��X�n�"�H�� ժO]o��4U�?�͖��@�z9A���ՕVk6h�"�?��w�nF�T}����VyQ,uqâ֨jΫ��a|�Ǥ��u52*�L!p��	���1Z�*9f��,ʆ���L꿼��f�۪�F��$X猾�]�6SY�P��V�����W;��1	8>ݗD��"�Bd(�f$��L�6� fߑ���7�$VP�/U�g[��~����F����r?ǒ��g�7�T�.y~�h�/۶�U����g�,�c9zp_��Ȩ�oqU�W6 *�Q��1L�E9D��޲jwHg�O�}��CA�r�$��!�v<Y�i1\����r�la���!'Qym�7��7P|~杞��	ߥ2͓g�GuxI�����8�~�[�xmQ�6G:��Ur�V���-x$&&��"JA���lV�aR?B���/
��P,��d��c�2��SC��]M-K�5�z�^F�eC2l���~�T3�+�g=n�z��1�3�V���g���Į����h	Nh֡�<�:�L�o���o-*� <r��Lhs�96K˙Q�WDM��q��W_K���j���m��(x��:8�BM���
`��)T�'2�w�
��̱XK�n�/��C��q�
�@s$�x�5�=�qf@vB���&. t�+� '�yU��,u�������5�d^��	�i��O�̣Uy�Q�5�&�f+O���V�"t���yR��sЅT�EX��B�c�O�^�L\�A�׵V~�ͭK�����y���pR���ս{�Ƴo=�D��V�.d�@b��o$�^�eX�,n.��ᆥ.����tD��%��UU�
�}V�5���C�V��Y��SG�m�NG�L���|�46�G�D9|���Jz5�J�S�y�s�T���uG��Y[�1-3�E�Q��U�	vv���M(R��m%�/2�Sě���E
��gA�bym�^� %����?b�䊳m�d�����f�b'��ö�v����Z!���^���I;7�wyxr7�a_�Xϰˁ�v�&�����(��wX�8弔VԿH
�@��k��#M @*m�����#3� ^�ɻA��ul]�.=��E�g�ֲ,��?&�w�����8)��Bɫ���¢�:*�!�Hv��0/� \� n��ӳ�N>}���Ԙ�쫄[B�d�><9�B/��A�ૄF4ۄy��%����w��(������EH��)�0�=O��s�1���J`�ci���Y%������`;9*{�|�Bn{����>=���� �L/��f��u�˰0���mT���qBd��7�'�Ma:&���Ϥ�'@"�a$��"�[��T�7U���tn�$|��s��#@�B�����F��l>��+s��c�͚�9M��l�5�RG3`��,Q�~f����]٧��wQ���&�j�o��o�C��Z���>����q7���"���o�ĺm�7�(�����s�c�r�O��B,�,���LAj"�q��j�sG��VN�60jӭ��H��!uT��3�#4"Bz�W%�s�7{��a�Z��±Mξ3w
Ld�V��`��?�O�_���t�8�����r�ju黖��t�R�3ρ���8�E$�Y��B7����r����������?�s�L������NS����c�g0P���h&�#�ސe���-�����$5'~&�%~�Qjq8*�R�=k��e	��> n��}�d���On��cA��h%�s����@1������O�&_�m�C�8��Sf��L��)�>�kqǓ�e�l�|`�d����J[�C<{���U���J�1	؇��>tw:9�6�;2�1���"�Yd�q�f@��A�c�pH�V��Y�X^+�%�M�.GaK���������mL�l@�&fE�Ap,-�V/u��%:�h�Ӭ�<'Z��	C< W��-����q 7"2`Q�˓���. nl���q��G��I��E���}o��$��f2�Y�x�W$r���Hn+�%��7r,�Dc	f]�c)�����FɭZ�Y������7�L"ͼ�6>�jn�ץ�2J:G�{�w"���[�	�� �+��F4�|���b/r�i+ۧ�8t�a�q�
�eC�d��o�P*���Ȱ�/�t�y8��������΂�NU�I�%�Q���LZYľ	�N6Ɯ̝pj�\��q�9,��8 ��u@/1��rW��1�A�!Q�(#n��m�r��~|lx�/�E4�n\���`z�S�R����F�L���.�=�G,~p�i���RÞ���vzPI�F8�!g��G�g6V*����ت�
�l�&������j-L���Gį�G�г,~HD�|����2��$QcI�������#m�qӲ�Ud�B�d���cvP��z!q�͒G��z4�QZ�(	�dF٢o2��Z�v��FI�G����������'A���~h�Nxz�1�kCm�#����9���{#�OQ��$�0�qC�t;Y�����^����1��z2���Y�k�eݱ�I��L`��	���ks]�Rs�E��n:�3�����żXf�2�S�Ǧ�l��n\�1Il� �$� ~��� �|W��--��o:�h���"���g�:c��$�F�f�x�| @ �uA�?@^bC�JΚk����r���d=�eu�0�}m���%�A��{�v��s�B꡵u�%ix�I�e�y:.�<�:��x<+�����A�GȀ�E���0�d������K|h�)�7l.��~�ՒI��)�{2��P�<� �����!���%.���-ۻ2a3h!�I�f9X|֫�:Qr+JU�����~˫_J5'(D�@��%�+V���u��*���E�xK��Q~LDҴ@V׏�R��{v�G��$�!����܏�����O�b����ο�&�\V$�ҤWn���TO��s%p�8x�!�|;�M��]W�WT��>�7�@Y��M�D��L
?l�7H���̨p`G�B����%�Yjũ��S?z�/����p���K��q���ZkIl�H�G���Sy��$R5���(�Y��� u�P9<L�n�C��K�;��K6%��άH��0�;��<n�H����/�<��B�'�-=X4�	:��뇲���׹ 4������|�#���Zʝ[�[�eO��J<s�i]��pf��̰��vڸ+'	�w��&w��@��^����6���\l�ea�μ�jp$�ǼB �H�I'��9������e������d�=M֜���[���S�A�:�ʻĢ}�
3�eX�Z���B����U&��DA	,q+���ɻv/3{���p؊��b����VwЅ���WH���1S��"B�[�+�L0epC�L�-P�X\>O��8V8�.j�����|�fM.�3h�V�d�f�K&����}�g��g^�]���]p<�y~�oùm��Y~����y<qV �g $J�h��l	���7�\��Lh��2B���&���~��<�3_euo��!ϣ3��]�TX���7գ����6�W��L	F�����OF>�7����
�v��'�{w�4�gc~,�/ܻ�㷜�(!x���?>=oTZ��/�3�Y�)`*�G�a\r� ����\��}�XJ���� c*�ey�G�ȥ7M��¬0�4gʊ_\�R����N$Fّǲ���F�Y���pr�o!"%�W�$
7<BoY�w��a){&��������ENW:7������8U�������~�T��Z=�P'��"ͻ�1��T��3>�c�F恖|���=82 �=�T�:HJ�N#fiۣ�����5 ��V�I�����?��_uql"���a�o7+C�ƽA�� ���`��Vj�%�m9˒��@��
�]c{�+�S7uY�H��t2ơX0�������=�N� �J�
�a�ذ?����g#�pl &J�K�V�{3�"2�h0����N�y�����Q7���X��_�`1N`d�	ז�i�_�:,�]�A$��f�.�SH���]փ���T&�Q[	�|�DF��D6_�`V�/k}���/_����"�)��YƱt����%y��]�\�����7f
o���AJ:=��S4��[/<�+�΋v&�k�.*��:��:K��~���>���+Ԉy�XV'�m�u{#���J҆�؞�JԼ�x��� ��v(sB���.$�=�r&� ��2�O�*�Y�DB���!p_Z<ay�Z��/~*w�q5�Õ�w�#�� �a�ť�M�Q`�z��֎U$��Ʊ�ѧ���}�{;�0WV�S�S�l�t0w�[�H�1D��4������]b�χ��l�)ޑ�X�)h�R�@�ض��v+�|Mj���c�r�22�2�pSھ͚ �"+@�]����(�&�r��#c�E���ڲ�fګr��e��P�1�X�lD!h�I�<.*���х<��we�F��쉡�|8X!BM;U���d�T� yN���S����`�j�{���FUE��"lU_~�0-���h������v%��U�8�1t�g3�>z�T�v��Cַ�vW9K���Y�u�� i����
���UC��"����h؋�N[4�
c�0�9Ⱦ�b�j�/{tC[�Zt��i�-�T� @��V�ج�+L��{k��7|I�5�!<��V������
'���]@�M*r<?qoh��C��R���gة��	��38)�9bso��ӥ9��Â�&�Q��ܣ�-�B����Xȼ�j[L��ҧ��@}ho
H��Hȋ��mp�*(I�w0;��]B���Z7Z��ic<CF�v3�H�0Ѫ�j�ֳ���x�D%$�RpŠ(uA,��ρ�BP�@����m�R,�6,�&�(�,����݀z�
��H�jYP��V�7|��熍pm^���V[l��jJLN�x%#���tW�\,^�S8v�:�m� �
�-�����0�b���:W�,1�����	�G��t>�̉1Wɭ���iFJ��?��gc_�������G�7�Yo�գ���9���/��RZ�ǲ�WV��?�O�}Q{a�67JK�:�h!D��[Lh/�b1ez�hR��6.@���Tߋ����O����l�AX�_��	SM���f���E��?	E@�:�Ŋx~�x�vz��l	�֪��0�����
��
	�ld���.�@8�'�<^����	�GnV��@���`���������)j+Lg���܋}��ˊ�fY�4�����[��<v����V��ZT���#�C��W��q
Z�w��N�X`�!Ql&���4{�܄��lD]�4�&�=C��.��#����89jL�IS.��x<耴���q�|��~�E�wY�凝ke���E�҈��n�
F�K��gj��g70 �	]3�֟��A��`ǐ`�.H>�&4���,��iYu�;�����w�=��+�������*Ē�!j�1؋P���K�S?8�v��=���a��9�j�����tE@�{�ݱp\�|��3{�KN�Agy
�вZ�q�:?@%�沭�T�I��F�~��ަ��p(�I��W����V�-K�B�0@$Þ�匞����N�5��	F���*3��tj��c��yVW��K��;51�r<�C-�1imԨ�OcC?)vMX�?��a75Ubjd440g6�_E����́)\>�;/NK����?��A���Xn��8+|"�X�b�����k񍤰~�Wogc�Cę~Z�8�7���=(��><IW+<cm�T�^�'~il�;;$Є?��~���Ua�
��h3��ߝ�\�'Ktt�Wn׮��
o,��b���d�e�b�Ab��F�>���D�p�9������X�M��U�I[)o'X�������{����I��E�fP�pF�Q[��[��W���&��r�\��c��cUj�X����,6�Hz0�j?)����8P����6:�@�XcĒ&4��y�C���╤�+���j8�wmA
b=߫f�@QP���W��FN&�sA�����l�Χ�7��a�ޯeH�ymR3d���&�Ʊ�W���f[O-r���d��JtP�C��-���zee� �f��-Ǩ�����*I�U%���p�V�R�/��,����p`���*	H��;���/֭rQH�h
��{�gu�Ap�6	�;���s�c�Ҥ�%CS��X�[���4%�d8",o�.�H?�oHQ�����/8�g�m�9D��3���p[��H�A�Gf�y�8 F��sFo��}�|���T�VJ�t�R;Nh����+8��o�zK��]�E$��F���U���ߡEI�R%z鐞/�'�34^�;�4
T� ψ���
R��3���m��҉D���E|UJ�5�!k�'g֥��Mx4�X �Y�ޤ���[*�gD�����bE�rx��ӓ�)@a<�e��7>�t��:p���Q�D!���:ږ1��v��+l|�Ѥ?I!w�� t:ص���Vf�N�	�Au��sT��-�>JX$n"-�uC���2�^Myφˮ�o��������c�;|����bH4�5�\ ����������������a�'��a��J4�ת�6�y<�˟���u˘�)L`�wU�7�]��7t[�Mv�N�f����_R\�*���S|�.�W����A����,t�G�b��|��sr���� ����&=�>�䳽���L�����`o���!y�ڰ,z�����,3�6����f ���2[t��A��X�T9
ҧ5��𴞄���Y��H��F9��*��]�A�L���r�����F�����h��+)�#�p-d/v�Ԉ��W��]C��ǋ�E��E�R��̑DDw+A���61�5��]R�6���5~�>�$�E�ǥ�@�-ީ�� ���"��r�+��uj��e"��:�9��F�z��*Pv �����;7K�ū�'�D �E� �H#��G�"��ؤӶp�WwG�L�����I��RB�:�7�x/�@YV�$�=Q�y$�_����ݶ,�<Zu|�N���L�UU���9�1��]�	��y})Y�qҤ��%J�+�Q	#� ���f��u:�s��9fjD���� :vm�4c̠��'�׬5*��J�����K��pS���\���'����9N�ʎA��v�����v�ɚ��S��� DR��Ӭ�S�������.��",]ˏ�w-֞:Eߐ�1�&=��]�R`�?���[p�Z>���6�����]*} -T���UR���Iǁt&��|+8�N�������)����m�9i�鳓���W�.�]$Z����}-Hqg{�H1��m�4P:�"�sO�E�h��0�����!�oK��N�p���$,�O&�3���9]V	���=7w�W<X��X\h#6��tc��������Z+"�[F�6�����j0���F� fI���`���A��t�s��_�,As^���K��C�w��3�'��t�Ϝ$����y,�mn� ��.���.��d��]���?Q��2���0�Q���p����b��V�Ug��-�h�?��߽Y�=�����n�\C����ɿH�v�4��nhv��߉�Q�%�J�[DU��ȋ�0�'N��@�~/G���Fқ����p�~���^(,S��8�i
�H����/��Z>�\x8!Z�����Yp@��pQ��oܫ��@����׏a����=P�%��{���xz�+�T�=׆��V��SCʝ8͊F-#*W�v���*�=h���}�s����mvb�ő�Ӈ7��G�r^p��2��M��g�|����f�e$��6P��Wu�ks0�8�e�%*����Y`��
ʧ���݃ڥK� H��6Lo�[�7�2�C�,�ł����
���"[��ȑ�j�eȫh�wo�×5�A�J΃<I�V��vY+�F6���G8}���3����a���]vq��
�@��l1mܙ_b�j����(�8 -�|_��e�>��`�3�0���8����Ȧ��(OX&ZnLh�S�V�V$��N��t�+,J;y_���jj�+��T�����%n# h@nG�	���l��r����ʹl\^V��6�o�$if#sp�'i�Z��2���m9�9�±s�T��P&-�h!K��yZ����M' �É뇕�����l
$�%9N��E_}`�'h���L�P�FS�2!S�$ٿ�R�؈B� �9t䫥Yz__��$C��ԕ`:q� \�-�ID߾ɼ���_
3���%ӧ���.)��@t���4��~_}9$�G�S�c��X�p������6`����A�m	�wR4���,]g����].�-'��1g0�����H�3Z���F�"N�q*&�
�����c��G�x�E�?�fc���	p����m����ޑg"IY�v?��O]��R������"n�y��yo��,�Th]5�$X�,�S#D��vm���s%:(:y��� �ׄ:�tf�^f1ne,�7&�`o�Ȳ���kVAD
G�k��n75ل��q9����ߪ�Y�K����<�}3��G�g^n,��0�\�wUY��T���*x�H�yGzA�R�.WE�o7��F!k�KY%�q�밺n'*���Wa����`�GOǟ{���Yw�� z��W�W"��{�;WQ3�y����'n:T4���c�t]��7�Z��xI �j:�9IC�)���!�赠�$��J�-%̥ �F(��Q���v����t����ګH�B@��6:��q���)�I�Mw��بL셚t��DV�G_�BZ��]�W��q�o.�ŭ#[����j����%���2p�i�g �N2��mܶ5%V�gK�l��?[�m��5�����N|�;�~�>TA��He�s��03��}�iU���{�UA�+;Eڝ[9��l�?�9�'#.[���,Ң��ی���2�������l&@rKb8��Y-U��� ������'"?+Os4�B�O��'	/�4������B�������{S�R��b2���otn#��!w���d���Wr.��~a�B�=!
*���Q���|K��2�_��nX��s�Jax�h|�\b_��F׊b�3Jh��Q ���h�.P����i�$B�*��U�Fo���T�BQ�L'U���%�\�d�'ә�9�S�$�L�}e����8J��ҽȷ��%A?M��wӏ�-J�;>9��gV���\��a ���3���cm������/��6��/)pz��3�j��*�#����I�L�R�ީ��{�������m*c�4����ߙ2��#�	M)��GE9�M�Z���d��
:G-VJ������ږ�ʟ���b@c��?���Y��ʉ7��^@Ĳ����Ab���_���M(w�f
�}��R9H'p�XB�f�I�ZM��´�"��EO�A����ч ����u晌��]� e��jG����w{�t�:���\l��>T��9uzl�"��i.��������-�o/ȁ೜���j��{*�k�O6}��{(,;*l�b| (��~g�:"�Ɋe��7���4\��˚8� ^��3��^�.�DO��ܠ%�zHE6��Ys�-%�Ј��ޢjҟI�.*�t��
N\ έ��u�,�
��į�8�1�:�l�V����h�H��QGS��o�¸w��Z'� � /�s���b�p��b��G�m�جXNzE9K�g��-��e��t>G���$O��:��j�� �,���Z��2�ϋC��y�[�꽸�e��a`� �og����):�k$��.ln���Ź�,�HU�(�mt=����[b��5���=�3��%/�p*��ƴF��\���� Ҡ���z��Oi�>���j$��
y�\��Y[�{���`3a���_9+��f�Z c"�"Z���{n�I���_�"�]5Y�|z���V�����Wh0����pÉ�w`�OI����piY�s��X�=�}���]jd�SK�w��Lf	͈1]�`��P�����'�mom�m'��Lvby���w8��|UPP>C���?%I��mԕYF	�Qq��%��PGz��Jc��rV�� bp}�'+���' �J��#�˶_u&�$o/�U�I��չ4{��F�}���J}7��:P�-���=ɼ��\�.'e��Jĭ"wz�;��'�ڽ|�a��_���f�5�O�zM�[8����Ev��:���t,3d��:�?XOP�|׊#JWXQ�v�U��B�H� m�	Lk����(,����S$̗9~ �PPN}� ?Ï̬5��?xr�-��ew2z�a%IF�]��ߴ���>��Q�h(>� bQz�7�u�����/����O�r�ir�;|�hB�*z���{,�%��p�	�_,s�4��(�߷q�om��#�x��=R!�ѩ���@�;V7X����j����i$D�%V��8E<j�6������x�%j+Pp����V�,��ny�(c��sPN2@�GGY$���Aov`��0b{*)]Wgޅg�;T�y���HpL�B�Wl�7��d�*R$F8p�YkH���f��ր�=����8�s�KAA^�Y��7����-0:.oVة�K9��M"-&����oh�[Q		kwd�!:�ʷ@5E�p��)1E��"E�J�DZ	,���C9�xOɸ�G�P���H�4mZA?Pg�;kG)�e���3\���1>�^n�{��S�h{��j�Ѽ�0(~��T%�h<�[eV�U�β�
�:c����R'��ͨ���Ĵ�?^a���cT
�󹁎��'��L�F����ʍBk�<�7|7ne��.YN��ѡnx4&7�+�'��U��Cks5�7t�)ж%�*�g?g�&�"k�������'�#���f\H��b��Qs�?O��\4f�:���O�i�u��1�Ĳ�돗�6��C*I���5rQ��+0a/UJo}HV����?�:�wL�b��o�kp�n/9Ü���~7rE�:���F?�1C҈'uWlT��}��$��Te����<�z���QEπ�pOh��k�yz
e��lJ�pH���F�*-q��J��M��z ��W�^ݤҀ 2�%�:�ۡxIS#�tm���Ջ��ҡ��H(�r�@ ��hu@U�7=B�b���7�6E�<�0۶}���6`9揁���躈|��<���R�".hoRx��]B��a!�v��v�CA썦��]3���"�?�L��n�ʞ�����̷H�t���u��&�����������R��]z��X�C�M7�.�S���F::wRu��!*��U�����t�M�W�̚!��j��܃�w����$��0ŏ����0\VI ��)"�Y���]� ��.U~�D�rȺ'@f���g��*r-�����˴��`S�px��Bf�>nn��y�|����Il��Zy	L'}?N�o)�oX�J=����\̜l��C43^;�?XԱ�V��Xr��aȋ�<"K-�S��=��|;����g}����}[S;˞�K�Rb>�6B��BU�k����9��7�Q�M�2�r[�5N�N�
��2����}�Q��5ԘǨ0�u�ʬd�c1A�T�7����	��%y)2D�U��H3}D�L��i&[���?�5_��I�۹����,��#�Ҟ��e��K����o+���jm3���Om� ����bEZ���?#hv: A��ŧ7��4o'D0��n�w�
SQ���Q{��w�m��ߦ���Vx��tTYmEʇ�Ok:`�PZe1ߋM
�%E���d�dS:��K�haL�ղA?S�9莡(�.�j���*	�t�r����r�Y�X"A#�0����Nv���~N�i�ru�����v,T	�M�"��/-�9F�oՓn���bi�_�n7֛��c�v�8Ӄ#.qc�&���t�;���Ӈ���� ��b�^���P��JE"��g�_�����$�0��w|޶�ѡ1�*�w�=*�D�{���j��IΆ���߳A�:Ƌ�Eg���]S`�����q�G�'ٲ*�m�U��0��O	��Oh�����*�_�1(�2�BJ+tZ�)�,��~�^�����lf�
 �ә����T,��N��f^]�˾ā�/� t����1�)�������k�*��X|���[���jv(��g�i�!6T ���O:r�m�����ek�3uEn���q��q��͙L��>:.f��,����[�.	t����?^���!��ޘȺ	�}�^�6���jԄm����ܘz֩��kt�p�L��blO�/�!��|��.����ޕ�����
����Oy�P�x���(dq�.E$�2z?YB����7�+�� Vên�9��d�`�n=t�� f�a�� ���YZ��ns�� #�k�̘aL�̋D��/��B����zFB�b���I|�x��0��^�W�/rׇ��xa�%o<+>����D���RV=�'k�籀���\�������^3>R�����e�e� Xm4��Q���,�R��&e-\r��d�`ʈ��=��4I�.=k�}�Wɐe�����"� �|֠zr�t���`J�SjӅ�[���2,+5�y��7
��7h��|��&�!	�/!w��	�D�F��ܤr
͗���7�	tdu@ĂJ���J�p�+s*�J�3B)#�����o�����%z��BG��.D��d�/��tr�8;� A~ ����b����,N9.�ב<���E�������lo�0#�����C����r��G�>��Jh�>�<�ބ6���������2sf�d�������U��i�z�ҵsEwҌ;��4_�sn�j���K+������7�<2�Sp���7�!��� a����Wk�~�g�&{�ln��c%����W�~f�}�"����ӞHXe�]1W�.���!�#�aAA.`��b��Y�'<ٴVF]�*�s߬����W��Z�ogO۔09��~4�ߋA�2��C#p'�_���8��F�����/�+��\
�p��s����鷘L ;�����c��[���3=�W�G��I�|8�Z
J8;�v E�3w�ܒ8T����مN�}�Q6C~�C�1��� 6�3��[W����G���o;Z�ܯ����F��D ?b�'�UkS_m����F">5?�n�X���'=��ee�'����-3X&E[G0��脇H�aR9��1��.�D�	�ʐU&������ڭ���[�XsX�2)�(�NT��/�������7M}�E�,�ꟍ��ڈ�qi��}9v(����bܩ1a��.�K�Pہ�`�\l�$c��}&!���j�qo�?%�.%v�&��ͼL���9��ƶ��o��q����ND�2w�A����g0ш_
���>`�ſ
Z
l~�к6�pl>�r�s�9\n.-��u�݃�x~��R��3��л��./���ΩP��QU7ij�6~Y��ۧ��A�~��XJ6L�Jrh��ޒ�W���b�A,�X��<x���n�Q,���S�3h�b���V���yl��[\�<Sw�������b�Ifb֥����k��y0�'%��\g$����Z�N#�$�qbe�l���\`0Q �9ʁ���`���\����F�!5�D#�2�l��4v�!ꚑ�	m݁H�1J2f�6� ���.R�
�
���e���n2u��C�c@��eE۴!w�l�V�ѕ`�.������<m�����j�)RJ���G�N�������ܿvr�[U�_"5ay�:��A �%�|��e;��O�ƌ�B��-�<+����F9۪���#R��D3��E���͜8�vU�x!�����o�3����բQ��j�ɏNi�nϩx�{m�B����;m�?6ڍ�m̑am�Y�������	���Tr�mʱ��A�.7�����$y Ѣ��x�Ha�"qd߰� ����g����D�Z��%e;�o{N����,\�و���`Ln��I�Q�~SUnh9�O�y�슼�zی�/jsM�NZx�|6�-t�	�Zl��z���j$�%�j��#�;6ؑ�cId�5���R^ 6��-��Q���NfAp�߆2�0JX�xT] �b;�#�-������Q�bU�B �G�jo@�ڟ'\��X/lF�L�bxe"��оᦜת�;8V�#�� '}@�(s,��fP�;ͺ�1V���hQg�;�zO�v#�T��vwOW�1u�a�Qx����3B�w)�u!J`��j��u�xqӚ�f^BK�3��,eV��P�Wäݩ���95;����e%v$��3�r3T\~�'&���ݒ��'}����K/8b>c�~�u ~�9��v<	�qͣ��_o3cg���,����[d�b0��Y���R�yJ��qPÄR�e^h��[O�[��灗�e�V�ZqXz ���d,�^)Y=���}w��*⥯�d)���^J��cO2@u��LKK�U"�Is�;R��ygEI*i(/��Iw�+��Gm���f��#��[����Hj����>��@�iO�Ì*�2!�ZGU>ʱ*_$�H��E.��K'RD+���#��V�Fq����3U��,iY��j��p����@�in �G'�IwU<�E����,^cW���b`Ç��G<��^�p�l�l=g����|�s?/|�W[��k&RE��)����r>P�`@�
�V!^b���y}�D 鸲�>�{�Q;&���^3֨)��E�n?�"6�8�mW�>����[.>~]���'c����A#�9����� a7ֺ�)�����.W(��8i�̿�}|��R1xl!����5��?���|�� )M�Gݶ}zݢI���MU�A\���������H�߉9���LȴC'�T�a�d��5�r��ӓ�x���E������6�N������7���`��B����Zxe��d:[���3T�غ[p��;R�1�'�C[Rf6�5R>/�C)+�ξ�M�uL2��s�8m=�D!Kr�������i�����^����u�jH�s����8��~��v&��s����2�� %�s�[�X-��[+ﱒl*ܶW��fi��*`U����MH��+�qx*Y8�= ��Q�Nc���z��\��7q�e�bt;�&�e�Q�5@�lfZ�\\a)�r��.�&�-p���7��Ә��SAN�5EC�c����7�l#���>���ʯcN���Y�_ ���k6�eM�?��K��o���ƣ���
B��N`�+GX����H�~��v��o�C��{v�Ri;<�k�3^�&�?1-����(v���"j��f�z%S�c��#��#��qz>��a��{��O��ѭ2�����з|�=�1��>��Jb�a�۵�|�`�c�S׋����vأP8]O��{y[�z(�䴦б�D=Ru��D��������&ˊrdIİ���֎{�$���.N�Vo
ǪKG�K�nC2n,w�b�+���oئ��U��r?!L��U�#��N�b �c7���1��=:o��)g��;�++m!Zʃp7������NN���B�ɛ�4{A�&��<5�\�CZ���EG�دC��v����=�;Ӕ!ᯑYS�*�O�5����'|��/�*���U\;�Y�R�:o�u���G�h^��5U���b�X�eJ��d�qF�(C����2�R���)dF}��u���q�jf*Y=��f�ӽP��~c��8))�
x�6�_ıs|�!dN����ɲ���:��$xD���>������;[�_�Y�l����-�Oz+I�r/R�Ў�<'�ىc2�4
�C9a԰?����@d��-<����3SA�z*�"�����������&F�([�lE�xq�g��t��[48쇂>_��J�I>I�ۨ�Io d8�4�WJp >�v���f�ئ�#�J�@��~�S�N��Iu�J�Á��|���8D�_c�y-�־�ɯ8�!�9�����H�?�y������
,�|�R��ؤЕT
I}ZpI��/'wޅ�o��.xTDmuX��(��!X�e���`0RJ.NU>`�O�,aO���`��Cӥ�(L`P+K���j�7�8������f
�j���B�Í�i�Ϥ�d���KPd�#FFV�Q�8(�1�D���=�I�&�B،nç���[�a�7��O��Ӆ���ti����Q������VT��ǜ`Sb���9v,���\�b��"�<r�~��Q1"ĩaȷ8O}�ʌ�&b�A�bҍƳQnӸ�E��>O��oZ�q�Д\��u�}��˞٤�'�i���7�Kn`%4��,xG\pMD��3��30k'K[	׫i��r�- ��F�R�|aq��G�''FQ	��ԴNr?w
�I8a ���T����mrc�L���\z+/qm��f���x���~�V�0�Ql��}��y��[m%��Y�:�ۇ�O�� ��SНP$Ԥ�',c�����8�<�*I_չ���pR���ƫ>��<������d��F*��/��t���pN�+��<�7�_-t��e5��:lPT3bl_�B�n��ü�wl@�����;qM�?e,m*^�
w(�~�)CX��mt�?�AlVkq�ض�Bw��׆v��{���s�W"��F��h�,��ש����n΄�B+[��*�ix��2�5%��U�O�=���]�~	8z�	92�G���R<<��
����M$� aL�+�q�t�uͨ��<�.~���ldR6�SB�C�P�����b8�e��a�"���4r��\L
$M�F�Ǡ*�-�>��m�h3��K���`����xx�	8�ͳ}���Of6�� 'H�f�J�綿�Q3R���#٩X�3��ﱆ�j��g���hf�-��vGSk�{�ߊT��c��9_"U��I����V��^�~J&����X��plA���=�����^h\��f�k�݂��|O~���
�b8�ىχi�(jk��Hr�+�C�W[�yz�c|�<{�""�{��&�&�lt��ICM��κ��OC �]C{HE�P����	Cu���/f��+7y6k�9e&A�$�w���uA��w��%�t�;�,U<<!�H���qS�~��9�ﶂts��܉��o�
vM`�w �)ǫ#��������u��V=o�o���������=@�G� �x^
��tmqr�|��;�/�`�W���>��l	$�q�����4Tf-x�vF|��Ak5�2�H?v��2��+��J�`�B�*W��?p��X��Nʫ�/+꺜��ny�p��t�x��t�@M�f��q�e����_(�7.��ǟ�;6hhwQ��J��æ���lQJ�I��x+)�Yҿ���&׺�`%^$I/%ʍ�m�mו{6Yo�����z���z�<P�@b��)�6bӶN���qZhd�� �t\\s��x#�q��_ߵ;w=!b��fL���*��LB�������c��3jH)��������D���\�\_�u�q�BD�%�'��eR�0�*IB\���$���̮i��Z2�TɃ&A2}F^���ӫ�u�=,�x�B?~sw�	�k���J��7q� W�����ή?$�i�H��ŞT���p����'�W����[�������q��/��I���i�j8Y���Ln�s��ͣ=�������1�Ƞ�Q1�G(/ /H�2
�v������`���J>$�Q��M:�Yf���l�j-��:ɧ/���I
��t>�{��PG|V<m�����		·�Х�l�/ў(�>�[��
�	M>Nv�zü�j.��e'%�˧�n�?m4#i��M*��1�n����׾p�5���V��ڄ�]��g���W���UK����Z�:�VFY�֢�>�D	Vm{�7A�Z�R{��~{�R��j�d4?�ǚ�C�L��w#vqYJ����U"���Mk��>����+:��q1��{	�/$�\���[w��qfWuECx↳��$5�����"(3o�@��31��g�ʫ�6��l� �q��պ'T;���P��h�����Qw�W�l'7�� �rc�x �_y���Z�y&;�����>��FޠtzDZv1�E�ɤ��J�A�D]A2��/�a��8e��OњW�r91��X����Co(�a_�Hw�m"�ȷt��u0U3 �Z�p9l����bf�ov��c����U�=�Ճ�L�ᗃ2�)T;��VVS.��dW������v*�&��>�8Ǜ���hf+/�4�gXװ��US�K&�Z�<�����wV��dJ�"�VHՁ�B*A-���W�DT�����N�Qb�67���9.}�;�Iq�[z;�$en�M�:�_��n>�xM��]^u�L���3��a�j�/�����-ky;D�t�#�;�_��QAQ|#��b�?���(,�z޴��^�>�$�=�GWka��F�I��OQ���e���)����{���y�C5�!�Ϯ�G��ZPFr����P�f��J��vxSꈯ�B��+�:�#�fE����`�J�J�4ĕf
t!lr1�"��(}�[�s �O���89���+L��k�X��^��3������ʢk��m�}P�*6*�>%t����������
s~0��]��I�A%.�Ny���œ\9��>�qB�Jm1,��>(�Օ��-�x/��B�>F���V�ـݷ��-�\����۬M�.��H�-�U������K\$����X[��O'� �Z��qrK�6L��Fȁ�@����P~�h�,��@e�R֍A\��|Mצ>�����L�s��S�!�<����r�Ol�+�MC��WM���~�	6P��`!�;A��4ҁ�����'��G�.� 1r��B(���ʚy�P*��n{�U�J�� {��$���j���Uq��{۩A���$DU�G�eyS�bF�֙	�O�(���7'� 
J��a��~�\ti�.����"��[f.��*n8��ɱQ�U�٘x��/f$�1�.�7@�@�IX<���u/���mqN?("Y�J|��(f�Dw7a�|K=w�pˢ�}��j��#7�v�aM��F^�5[^U�L_�1�o��|���3'����IM��e9!3A�<j��X�,YwGo(�b=�"��[c����Wf5Y2�z�R��&���V�`��L������6�ޥ1�W.g[�!:c��R?�όT�캎�BgN�V �b*bJ1� ��܁�؊���aŻA����"��T����7��S�+�w���ﾧ������ۍzUj����q
����U�j`�cB�ƺ�}��_k
��Z vY��jV���R�@:�aᧃu��MJ+����a5�o��!q����S���\@T�
��{x.P�����p�iķ�!o'�e����,�)�tA�r�y3eF�.@��=�`�_����n�����;��a�;��(}J]=���'s�3*���I[��S1�+A񞇧ⵙ�pN��]$9���^��i�esa=Я�DR/��l:��J(�m�n��mX�O��N��a{+A���ө1J��1ϮNDju�ZrD���	����NX�6?��E}�_��2+�)�����"K4�䚙m����׼N,���'	m����T[	�sT����F)�c+�M=ၰ
���*���7������1#�|�?�̮��NV�݊9]��Z���g��ܽk5(�K�Gh���͗<,�1wW�i���<��v�3�G���k&{�w��y9�"�1�s譻�p�S~0_�݄��d�!�&�^�3����LE�1�H7�1�)}M�8�G�.�b�ia� �ű�uP�n�$r!S�$�t;~��E+�Mk)�Q�غ��/E9���l]E���uD$a�')Ӊ9�)�!�?��ȯ�zs��%:I����g��rL�6�e��8�M�)B����%n��>A��{���::m��o{!��J�3O�m��3�ò^���j���G7;��!���8O0���s�2f�!qSzX#b�5?S9�*�B�x�'#���-R������E�<}����9��O$��P�u펽 ����:Q!���\ᖌ��ms~���$�W3BU����T�_*�������++�c�S�Q-�D.Q@�T�q��ض;�3
����c����HZYaw����
�EϦJ�S�\�B�s�g��-e�QKk�B�S
z��#+T9�Jj������̆%���e1�@���W�֠����C1��z��8-O����X�S��'�� -�g�(@��3��(`�[Uw a�d�I�z��ux��qbm2������J���b=�u� ��l��(�ԁ�P���)}�C+�ʔ�߶�h􌤯Y���X�2g�wl��8�}@�U�D-�J��[{(iKՍ,��ֱ�����r
W��\����'۲8����]CN�>�}���cYR��I,!
�hv�V�L��1&��]�#2��U(�z ���E��G65��'&���a��o��N]� � 藏�q�h=|~4�#ۍ�a��m�"5eX}K8ݳ2�V����<�
�t9���x��V ��KU���xL�M0�pLW60����GNv�o���עz�m7�ŀII�C��X9BZnE�u4pR�p�Uؒ��$�f�m��Ä�<u�Y �D �j���'Y]z�׏X;F��G� Ƀ��đCL1�T�5�P�\9	��Hh}/h�=�L�"�%����وxk��D\+^Ր[��cܷ��1�<��A7&���8���	TC�=�vB����C�ة-3��Z�D#!w�{�������G '���N4B���U�&�/���R*��Z�G@�Z�}fQ5�ײ+#5[QH��p�����>��}D�E��ַTO1F�V��d"#s�����%�-\�{W�������֜��2�����p��oX�ͱ){މIAԃ�xވY�{��v�[ʣ�6Q��_�&�����d�"�W��Z*Xׯ,_���phY����z mfHt�a3�����#���*~
C�0����w[0�|eϭ��;��i�R��Ekq�2�i{�@�̦)��a�l��hEj,�9H�2�ʛ�E>.� �M��Ͼ�}��I�5���W:o9��oj�>����ʲ@�<w\@IB�+~烂L�[oX�.˕����� Z�Ʊ4���/��9}<�w-����L0d�!�W�l�Y]�j��H�_�5�ֿZN&����C�>�m\L6A{��`/b=�� �������l�j> ��E�-Y���V���t����A��`��fW��t�rϷ�7p��� �E��h�
�c�X<p�+����!TJ`�KRJ�ygݿP6�5Dk8������ϻ�M���>�9��ۿ	��:��,!�d\�IA|�&�:�vq>CH���&��� Vk����YL������)�k���X=f��vF��>�"z��$�ۯ���^܎�~�
aA��N:�����U8�OQ����_$��^]�0
?Ot�Gm򓡣�7@%Q�a%�A�ԁ����l�ӫw�戥��=1r4?>/V:�,T�Ǧ��rc}��RPg��;KW �?����dm^�i�&�#�>E���f�Ζ�p~�����f��6�+�n�X��6��2������|7�A��%��ޖ��n�5��-�ԺaxE�c�w5���^��
��5����Ƀ���҆�|'2N�#�Hۋ!.�vڠ���=��g�A��=CKG6'�М���vA�ک"�sެ{L��~1��R����+
V/���DOkf��Z��|f��I��v�S�#U��>�}HQsH��E.�`/;��t��j�_X����*�����e� X���Mצ?�h�g���S�k�|Y��/���<-��!�ۥ}ϣO!:��i��9��
��Rr2ry�n�+b|��4j�j�.R�����8W��p�E�}+M�K��6p�i,Ə*�|�u��;��іa۾e�?��\�u	V�mR�sr�mp_���5o��`�f�����u�]UI�y4��c&wo�3{H# ��'A�([� %��.����zV}'[|���R��tҍ�"5}F�+�\���΃�1`!�.m"�z��p��Ɨ��:�Ѫ�W�M���8@9C��/��Q�r�%�uE��g|��w��� 	x�k.���_�1��&w%���En J��~/U�<j �i����B�r��u!�N�a·g��7".QK�gt�q�4����~>�&���KJ�ɱ,(S�ꁬ����W���,����7A��5�������g8@���BBf;���_��	?_;}]��Q�	�3m����)JZT�R��~<J���]&�|�����4�W�7�� pV�aJ\�^A#�� ��O���6�蝰����J;��9�. ��KJ��Z�ϝ9�"m�]��{}&�^��AA��I��ȧv_�=�_H�݋`_��R:�>,)�2�J,4���w&�#S�-ԠD�*�����®�6m<���p���0C�ѻ7����p��{5wq�=cX���>i>�h!G{��.�0k&���4 8����|�WG���G��0Z���{p/�L�WQ���t��K-j�U�'es#�-�GF�G�(�
ET���iE9k��%
��#λ����N�������s5�qш%�k���4�v��w�iM�;�8����{��"4�������N�
%�r�T��o)�8��I h�2\�y�Jp���]@�B��%����_���/e@VU&�ɀ�K�q�p��#)B��9	����~�����cIX��
'��j� �H�^�+SL�6�D8*�ҍz��pni�"��9�V���\׍+����'gǛ�;~(*��96�����{�a��~�G����m�Z�\�_;�D�e˼�~U�aɨ��I�o���J���Da6iV��6��,�U�2�ԌAr��CLcq�� J����l�>~��݌����7@R{�|= �q���c�ă�z@v�> ׸�[�HLب�k�v*�b�_�N�(���?W]�>-:!�~.}��_qoG�ߡ���Km��=�u�� '�_�t��s��ou4SE���g�$�&�Tk�y=c��n÷YsVRB���q���;��}쉀�b��� lN���i��,qP��p8�bŝ	x����A�Y�pf��d��(}td�s��D��Z�7�#�{�c��`{��q�n[�~�]�`���:��_�%S";U�u�#�u%��,�Ǧ���k�\zɱ��N=Eh0ɲ齃� �d��|�rf�Ҟ�͙K䲦 v�:�(� ��k��X��0���*I���|�8d���U���J	V��W��6�eR��A��e;�E.L�닖���)�;���^�f�ً����;��o�D/���ħ�C��o�����>�'�������k�)f�ʦ �\�s?��_�du�N�xv�f�T���_���
h�x�мC�⑵��2�Y��l��p��a"��3��_��u3-2gf �`"�_H �)Z5v '�L=�%5��
I����ڂ������T�C��8^R#_~��C�9�jN�qUǁ*�2�L�T��|ࣦx�,�����+jk��w������g�`(��?j�F�e:�����ʮ�(c����?kH?�^.Z�ؘ�v)�or�f�=I�i��<�Gf)pP����9{mw���V�ٺN��zFO�p�DM������ƽ/�i{�X�s�B��15y���k��V� ��*�=qݭ7���4��sֳv
�	�	�غ,�v,��ci�$�:��a����K��|�iK��)Sÿ��.�&���▽dw��M9���N��DFWӆ�f�͙ Ȅ�����6��Ēf(<�Z*G�ZU:�h:�6~;'�|q��˗��)���C������Yh�u�����u,h�b�O�&8Lz�t~����N�!J�ŗ2��f�v`�%w>�̟4Θ>#%���/�x�R<��:
��?�N�2E�����J׽��?�P���FҦ
~k�ƧK���w�!0.�+<�qkm���������p��#��5#� �X�m��*�Pe�E��K�}5�+���7�S��f�!,��z�(���j� =�y�2T�)�ʳ�H&����`�k�`@+��uSQF'��E��q��r�c���/3�oo���[P�6V֞�2�I��W0�rL�(qe,���!]��Y�ŗ#^/ዼtb��v
0�_���9<�fZV'ŎE<�^ڟZ횶
�Χ�i~��.]�H����!��ԕ"��L4��ib�
�gTM-�:2t9���`�����?�!1� 62��P{��`a�����J�<�1���F�U��WN���՞�=_�`z�nA7P̠뱗_��>K9:�=C�>L�k�s`6��e����W�Y9d��Hઉ?�zj�=�v��P.A��b��2�>�?��-�O�%�8Q���l܋%v�x�;���8PM���qk90ڥ�n�~�a�f?uU Z~�S��%E���Ĉ�B��s2 	��p=�k(yytx~ p0{����2ݞփ|���Zg$.�������sExj��@Y�$0�!a��_H">����tT,���w�@�,V޾ �����*�1Irʩ���h�$x�+'����h���	�a fMіn?ya�@4�D�a�`d5�"���(���kv��<m�&��w充���XO�in\��ꇆ�JTcZӔ�}��0$�Kx��0��A����ϒ���2��Cg@��5�x���޽�p��S߫�SW�ϸ�<��L��[�?�?�@v�w���w:�{43�`:�Ř���B�S̖9l��T� �ӹZ~[v�0��=��h�B�y6�}��|�&f�:�[��e` -����{W;��	�9,�xC�ͽ��<ԅ81&��A���_W@T�;���5	3�����L�^��̯Z�Pt�Wd�-������R:��FL��~(>��脴�L�f�ӥ�J��}(�Nэ����Y��q�?i�ck�5������O��{QB�V�w(?����ҒH͸�:\�#��e����XŅ}^�k�<��O�"�5�9��#�F�Ť���A�	��~��E�2dB~�O�JZd98%�i����~��2K�~k#�����w��ҥK��6��ۛ��3�f�| ����	|��QZC�W����ti� D{�u��tAh�fg9$k��,$ЏA(k��ǲg�%~�]����(����M�ynvR���^hڨ���yfC�(��A2�ǽ�b#M�W��RDX�5|�M�$Q=����{cE��^��M1B��t3
6fm��\�B/�#�~�q��}r+L�0%#r	�sZ�,�k�(�e����̑�~��H��!�"�⫘�-� �?�	{�C	��LW*�uI��ȝL��%�b+�SX�V����E�	E�+D�`�	=���L�\B�Zr�z��e {�@�jf���[�n\%�z@�����/����϶V�Gt�R��J��/�����\Kz�fU]r E�O+�����+�>c5d5�?�4!텄r�Z���}ǏDa�ם��-�u�y�z��ӀW#�A���^N5�׏�����M�%���+ۿ?ʢ���먅ǖ��B!K\R
,%�$�yS+��r��KN����Z�����"��M�s͉����"�At�w�X!i�ʹ��9Ή��(�k5«F0]��~k���ʋ�+������sh��s�Q�N�h�W��_-'Dtx�;tb��b�po�cS���m?���ør>��_��\'	�5thz�E��I���h��;�Q]$z�6^�M��E�Hf��-�7�w�#|������bg���v���@]�b4+���s3�(�c�kؾ��*S���\�͉�f1+oZ�1�yg��@���3cy��� ܜh��Ŧ�T���@q� �ɒT��]�XA�_�@���Gi�MI�+����S��p�1GŖ��+v���\҂�qc^&�u� 3;�и1`����G��^0�@�j9!���ҟ�u14H�;<I:��ݮ׬����8�%�&L�k���Y�O\�a��_���J��Qz���=�6&E@H/&�Nդw���.Y<����"M 0L��u����N�5p&��J�����t��YIy���n���ƍc�QdQ��h>�C�E��S�hf�#�n-���3��D�Z-���|���!�5sg|͠fj�R��9�)ۣ��Vcɗ?�-��T�ȍ�����t-��oS�2������cEtc0L�(�7�5 �rǺk/�16_EKL^����՜Y�	�&��	��V�t��6�a�����(�]h����G�$���U���^lUr�U�'$�JF�׵����,�l"w�Mfmx�x��������Z��Ѧ���K�5�����'��y��&0"�|p2c`�T��F+����ha����3����냛e�G{�.ȇtP6�%嚒J���͏g�F�D����G�c���V�����������vBS
�q�r�m.��Br�Ӽ�<����@�&��kh��P��=�a�+`�Q;�2�B	S-���7ʣ�Kɔ�22тT	O�䕂\>U��H6���Ć����"㤇ک�Av�n|;��O�c�sY��X��a���$����O�;�'N��𧓩����pyk��ʩ��ۖ�t@}���80N�M)<��:A��d$��éGB����AVd��'1�X��}#���8w��B<1�X�nv�*J�Rֻӏ!4|{�*J0�7�v���i�^F����
���u�/܊�ʰ�+7d2[6��Z_u����z4
��[�Z^��:LwB-� ��9�sOv���"�Dl����\�L�����GS�2["K���b���s}jF���D�E��*�.��Dt�����ׂ����ͥ�5!���]C�w��]b���X¯,��֡_Pz�'
[�����M�&1�ۧu�2̋U�����Rw�Bn�ed����°��{�t���)(�ɞ�D��`����d��=�4f--1E}��I�tӈ*Þ%��G���It'�K.N�>]>VkW^��(|}M0	�@����c�s��(�.��¦�A����U�bzF[�QkҀ9�@pd�'���D�I����q�;��N���f]u�9��A�k	#s�ט]/�����<n��/�K���2���g���t�����ir��a�����]�.)
/@a�*�U[$dW!V8��)=�=�P���� 粉B
��tבw>�X�<z����b%(����B<S��I���������~���Z6'���>�[y�}hH݄�C��~	,[�]�(�Xu6�d��� A]�>�k�����Ş�jRHO�F�Nq��&�
�b��EnY����]p��RK�1{.O����p���W��{�O�A��x������>M�%hT����h&2=-�3Z�k�(�by�m�l�Ϙ4��Tc���)��"���?(�N�1�˄X���֞�a�
���@��-"�9��MpE����)W#���a���zt ��
���_<K(�(�]�>���3�H�Z�'w�Z(@��b��/!?��Ɍc~�$]���i���,� ]�R0�2A���y�@Gy��N.<�I�G]�����5-�co���jl��8n�%��@e��j{����sȯ.���.Ђ��ln�#�4�%�%���ӵ��*]�L�Hv�=CJ�_�U�|�V����\(�E�+�:>�V%Z�5M��9m��u݄�� (S�Ea"�wcg���?//��|��I���D���Ofs��u�/��-c%	�9%J�]<���̎�my_~f>Ma��4�Y*�����5�/���FR���uA��N''H��2ɲ1əV�T��6�=����kq�(2��9���J�ύ=d�f�L�G���?���+d� ǝ�&7N-��i �ґc�sߡ"�b]6�m5�A����l��ӯXu�-+�#��We`�ơH��6��db��t@#R��Z=֯����r��1��OX�R���h�0����.�0��N��^�}����Z�I'�N�x�UK�7���p^���g��=�!ǐQ!��A���7�]W��#ˌq�����_f����_m��VpM�*�hp	��Pu:��7Mh�cK\�<�4�!�2�3:lh�!A%o�[9�k�P샒���k>s��sTU��]=���F(���D˨�͈l����x�0Z���瞴w�2R��ߦ?�^�;�n��;g.�xB�\8��*(mL��ˑv�T9Ǳ�q3f��@�Ɔ,�����)o��/
�&H��Z����L�D3<��?��Hs���p�k��]Ѿ��;����{��ik?!Q}����`$�0�����g�6�Ѡ�l�J�gg������9�}��T�cu0��<~?�Հ�S
�(�%�{k�wD4��p"�J��^�2�S�R�+N�;�W=��M��0�(�6Թ/7�sQ��U���`��I��2�.�i< m�ߔ��(9��� ��at,s[ G%�0 l�6�p	?�Z�N�̩=�����Fn� J�Q�u^�@�?�&(�K�_9ڦ��9��s%�<�#a|D��� |���kdj�m�4�O��^�fŚ�ݩ��$�轍p#�sM0��C~���<y��VW��5B�H
���+�^�t���30���g��&�!]���|�D(�!%\���g����*F��I�s�$���ƒsj��^�(�&t$Hؽ�x��'+�v��&��52N��)rX�U�5��Z��VY��=�m�x�7�n>�O� �$Dp�]���&���Xk��3�i6R-�Ϛd�ר(���Tx_\5�kC���� !NEʳ_J���!�T�[2>�WPʏ� �����t\��wA�s�4�m�Z�:M��3�(����b�����#�:�5��]�"�6�.u����>���!�6j�~H�f�qi��u��,�W�~x�B�,�β4>���>Ur1��(,앗��e�|:񜈵�X�)��iOl������+��x$/� 	=�ҾE�
u0CF��v�SN>zG�˞h���B�-�9/-�
���Yk�N�^7�|4'�����bT�Q��t����m^�t��w�f�p����Į���֞��ǫ�I'e�����9�'����p>��2�Aʞ�{�;lƹ̱Y�~����"-g�}
�K�����~U�o.&�p�ei��t�_����������gx�Q��k��yA�E,���E�)�/��r('O~��г<춦�!,�y��^6S:���|;��M�6�C�!�ڰ�!R�2�/]Tۜ�႖0ֺ��CCd�9o	��:�����e�F�@1����w�6��c���JA�3Y����m�(�4z��e�s-qP��\�n��l���#?t
�W�����)-B�5"dR�-\��ƂB�Q�J�K��.\6��k�zc�eb�'�2�#����N1���$�r[)���B�R��L'2�,Dޘ��h/���Z�mN����s=�*�}4�Mz��1~x��[,Aba5p�Z<@$����gx���z��ٙ@1�����np��* ��A�ώ�����}�{�[�>�T��'4�4a�i�a%�#��gIĜ�N;Ǟ�]c�x!ag�9fR�ӡً��y��H$��C�%mP3�"�%��c�hE0���f21s��7��0���0��[a�@K���T̯<�̇�&~Z��htd`�a0�R��؋�&��K+���ן���b�2��||%��:�����e�ir6{2Ыu���7A3�X�t�*�)��iQ@�t''B��e]/7����Y�L�m�m�����b��l�&����{�>�b�m��a@�g�H��7��Se���Cb��`�`Cg���
��e��eqN���	�}<͉�e�ьe`Ki3�8F'�dP�+{v��<
�Q���H��U~}�#�s*׀�R/bߡ����=쯱7�/���ea�@�5�"ńh[2b�� .m��:E�V��=�Ku20�C�B�G���S^q����՞�+/�, �n�ͽ�M�/Pz��)��1<,�T6iV �x��K�N��.�������{u��CD0���2'�12c�|�DaqY��[�ڱN�З6�Nӆ{3ɤ�REB�z%K;&�4�%����n��$Hf+���ɽ��`c�6�\xr�Ilʿ�Lї�Fo���-����@j���͉�i��劓�3ԡ��	QuS����$��Ь��%�T:xчAK�=H@�0�H5�\-B��Ս"Ǵ�/��P��Q�/�`��?���I�z{�$g���B����g�"��^`�2/�Z}>A�i�������x��ƃ���>�����pi�?���ԓ�/>�ѽ,�&��K�ܙ�g�����*�jPJ�}F�5M{�J�=p�J�y�ɤ�o����?b�ބ䜗5O|rPF�-�*wn��Ja��!o.cy'5~t��is�PbxD����� [	�1�����*#�Z@����y��zh%g�"�s��%t�z�]򇧝 J׌����.`��:�@{*5�X�^m�+
:qvq[�p\+0� ���P�@���w����ͻ�Yt�Π���h�c:��x��b��jEɅ���#�_�I5ϟ=� �o%���5Y౷�ٺ�\h9K5;���t��Y��rO2�
�5��2�`I+j=VB��`h�Bt���e���C�s^V�k��J�}=���B�e�!�r���a��f�o�k��N�ڹU���Iɭ��!��#M2.�!�(��,=(l ���U/��}���t�tE�i�a|�l��l}��DW����N�P	n�77�]��RT�c�<�
2��}q2���8~}9��ܘ��?OsF8�b����sO��r���#�>�OS�/�9��RD��A{s�����Ɣ�WG b���?��I�ߚeh��Z��h�L�ob8����IāH��|��4���n��@��Fϭ�k`4�v/�i6�מw��7T�Z�md�0˱N^�wM1����_z1(�ny��pqŹ�1T` �C~G0K���4p�۩E.׌
�d�bW;b �ٷ�r�Q-�G���	X@��ѱ�@�He����U���ͶMJ�;q;h5��xYt�i�p�u]'��Əmt��ctf�3��Vh{�&{~,�arV�i�/���}%�����&�.{��!��v�f��n�2�J�����[.�L���/r����o�5�P*]��:>��\��ɪ�졒e��N�(j��Pv�f%05��v6�:�=3���nD�2�YB�"��7l�{;w�����8��<�6��%5yTgd�*wц(V�X�q~�6���������v@��&�ŸZ���mi�����]�7����5�G���*��;��KOݞj52�gHy����]�C�ӑ���ߐ�)��C �.*���3(��ўuZ��U���~Qs��ޤ�������$k@.3Q��+���F�ji����P[��ߏ�p�
Nab��,�t��kxB��R�1]�+B�1Sƚ�ʪ�{������edR�w�I�\H&������S�kE�w��_�|�Y{�F�.Mk����z�U����GN/9��SƤ�'�/������PL�V���$�f���q�M�ߓ�:�h�@�;����g�^�b��La��]�Ҝぶk8���Gp��+8l/����z������e]�R9{�GcЫ�qm"��c�
������Й�B�(R�$S�k�'��G#�`[G�1W}��(��$Qa��f����e4�}�J�C ��d�__^Ǥ�GX'�+8��h�i-��E
���^��D�9W�=0����b����(�v�]d��ݛEHᣠX�H����K�x�֚ۤ�8fK4� ý��b.�g]���Kt�1��F��~�nq{ĵ�Wvy:FKw��q���1�@�}�#5"dN�QwѱPnd���G=Ϟ�o���1��:�#�c��E��<ڷ9��/�B��m6+�a,��h�;_G��U��Z����z�A��!'qm���Evȋmg62=�����A���i� �ý���L�V�1oP�|I�1e��_�3#�U���r>��ejHs��l�1��(2�����z����f���-�UU���.�&*��&:��?��e�qrx�|wc��v��{R����Aa	d�#��*m� K��,(��@�q�w����8���"�G�[b��ێ���r!�JQPؿ�M�<�����l0��|s����:��W���Y���>{���E��5�B����N�h�}�C��W�ZYM.�'4r{2e��0j��6r8�
��/�\���\�:�����L-��c��U����3(����w�$��)�(����h ���~�{�Hv�3������� SN�����S�?�W4'��>9xM�����ŇJ1^_���$����ԋ�[5��P2{���"���ۃj�O�V��v,N��a�}�xӸi��q@_��2ȓɯ�y�lEvq@D���Uĵ�b���C�ʀ��ĢMkat�7g��H��ڐ��w�wF'�Z��d��H��b�ӮHu��"��w���L^�m�CX��h�����d���_�U��D��fg�HI���u�+b���R���A�5�.�8/gJy�߿�eU�����B��.�e�=+����/O�m��NRը�!}\�>ض�ڗ�n�4�g�(�Ռw�П���10��!�ïFQ21
al�, ,���oG�+�Z������7̍�*�+P��޾���N�<'4�%�
8
sOjȮ`�2@�����[WM��B��@kOK?p)���*l1�`��y��Z .��Y�q�Bs�v�[0sҼ|����N��`��FA��Gl$��d� a>gE,T���:��|���=? �BGhj� �I�m=QW$[$���e���#��_��T�E6A��i��u<@aUA�\��<�q�ٴN�`��#R���e_����݇�9��D��@��(\�L|�z̪ƏU���z��kC��!�h71Q��f	�j{�J�2HY���x>G	����A+�������0��O���߶�<.��+kqy,c�9�9�b^۲��ǣ�ϯ��S�r�欣P�� Ʀ&�a������~$/S߰G���m���SS����J9�p�a�I̅�SK�R���U��u�� �[>���"�}*��º`�Y����ݶS�'��(T�	���4�TZ����T���_2��,o�i<�6st�b;�3�'@ ���!�i�����/��O?���K�>C,�9%��L"��=��f@�xb|���۽l��Q `���r���]A�3ήM�,a�!�� �ם�&���T�'��8ʍ4-���At���1y\j�T��}s�1
��G���z��8;-PT�2�_XbF_V�~�w�_�n�(y>��\�Z�đf/���>{Χ>1�	_6D����2"�����d� ��X=�&�y�\�Z�H�9�M��Ye��/��q��R�e���"����qu��"��2�$ٱg!�&�3��VbĊ�� ����8�$�T�c9�J�/�B-�R�HI���%@ P�J�U'�����Ļ�S"����/�aSm$	6�����*��~Z����,I؝8\��k�niJ�
�x`�TTEKƹ���7��sE{�G�����T�	�x�Ŏ�!S�;�e���3�L�m�I��n VP��([l�1��}F��Ko���TjEM7�����"ԝ*�l$��9b*��  ����e�Fo5�D������T�nӀ��'�	�!W����?�?_)!�iW���/��w悂��������cW�i���}Y��eS��L�V^E�\.�ƭ���h���U��fP�ы�!45�jJ�p���>q���bޜ�4���,���0�~�W��@E��w����j���1��~��Ao2H�[�.(w��El�A�$���b>ai�4h�;���Λ�~Zg��bK�Y�����w)1�����iV�Fcp
�Y�#�讹7�I��V��T�+�>ܦ�A�N�����q��������)�8�'�zI! k��+H�9��
�ס`��k7�ɑ�	��,1�.�SRF���zf�/���OG�V�i�ȃu�1���ߏgG7Xʁ4�/�,V*j�� ����������>Uh{�<�
�T��=7��u������D�?���ζ7�N��.!����$gn��d�������Q���;jIR��c\���Q�	��rXW������&]��3��~}-��1
�\��X�q9�z�}�X|�֭mc�rt_���u9�)O<Qy9��a��<�b�p�p�z\0�{���
��
�C�C�Ö)
��y*a��xW�Γ.�bHW$��A#�R�^�f�����ȩ�� �Pw��u����Hz���qJ8���%�OÅ�~�1S����Caʸ��*���n�I��5��v���i	���kO��o�����Ɯы����L��{z�@"�q��)�✃��FrdC)^�;:a���|_W�rf��pGl%!������$~9�O��C��ɫ�ZC;a������!E�a/�����ضK��>��N��pMq���pͼ�w'��K���/	�Ĉ#��]�����5H��s`�2�qJ� +�7h���ޝbP���w����8��T�҂a2~���W���=)|`'�[�Đ��I)]:,�+��0g���[�3�f����[��	����1�?�ķF���✞K�<GG�gL��X�o��G-��<�x�8%cS5_r	�4�F*�[|�_�d
��ndIڶ<'��s�Y �2�|B���|w���ɼ+iR���������w<�@�ר$�7&M��C֘?	1XZ�vTD���j+�d���Ryъ�o�O.3 ��0�^��&Y���8��f/��5b�	A
�&jxE�!�|C��=D�;�������O%p�!��]GFp1�u�y�������f�\�K��Ύ%޽�m��]��6�Pt8W�S`����Ke}�U^UZ�v�����- %J߽\(5v��,N�L���z�@K��{C�1`��p_�xD�9�y8Hb��q���;u�aq��'�$�m�Qz*�E13��c@�B){�������:uX!e5�0m�%Ɛ�k�U-Ɛ.�E�+O���Q�.��;���������!T��r���������D�����"��e��	m	�ݫ�u�ϔ��S�:��I��+�fϷm,9�UT���g@X&1a0�{�< 肻"�u�~w��uۅ$���_�����t�����	�J�(d�5L��:�<7�
�^��e�5�)��
�\�b�x5�S� ���&�$	���~h��n��|������W��KG���F�̺0�(sЕbVF��l�K�/W<r���%u�S[B��6�x�@��[��N�a��:�ي$D� hv4w�NC-�w#d�8�A%;#\���羠7ړ��{SP�.,��A<W0${�A��b!�� �DK����d3X�KbƂ.��	Z�" ���:� ?@�6���(Q+6�S6����h�O��w;G���J���o��M�Fع!�_�w8�"�����P¤�Z �vo�G�-���V��h��1q�i*�#��H�6hP4��rqN���T<���6 z�JJ6Ә��f6i���4����#���t#���:�?��V�y���)3+,9�Y��f�$:^J�&J�}��Xi��޾Z}�9!�{Ϝ�k�5E�h��G���X�?T������/m�;������D4$@�ELD�c$�C��RIbG|5���}��O��LYD��\��) 
c�#�c����$�[�@�ף�t��{��b���=�}g�%�s�H��emm��m�'�h��[D�����y�ip�/��X�JKr���	2+��>;�꤁�>����� �ϒR����<\��y(�0�(����뗃�0�0�5Y�D���RM" Y���_� �06�ŏ
����U�(�����t��VE(�G_'�oS�R�i-�5�z����0�pS��[)!#�a,/��Б˕�Tǝ��n�^� ��[�(�D��� �.?�F����B]
����9*�Qw��imc��ۦrVtc��qE�_��K_�(�t
~3�C��5|��:k6ubI�����"��S���R�HT($����MtǛ5�a�ɪ�CѰ��T*�x��e�qQ�쎐5?Wfg��h]R�zԱYu�= �@\y��7d�S�KE5�H4? i?k)��!h�,/���PoF��܏���s���ບ�2Y�� 9��ib���G+T(��k0�B� ��rh}P? ��s�3��-��虒�-���S,��4�d��P<l:�����o���5{�����g�\	j'�?�ږoke�z=�t�ɕVǱ4�V�
�u�$�(e�=��m{����n+��տ����z�)|�����ҧ��icʈ���ShT�'�D����-��p7�R���$gR�k�L5�W��I�{&�tuY41�{@������p+��[��ȫ���;�X�u_�/R�rEt�5��ǃ}-О
���2Oa�介`3_hM�m.���1)A�|V�J���Pٲ��o�e�-.�2�m���s��6�Ͱ)�o�~���Ӆ&�jH�Z�Z�^���D4�L�h�U"[2��f&Z�k�<�P�Kכ�L v�E��sn�ۥ����EG�MPЬ�[�}���>9�"�J���1*:�>�#�EՖ�B�b�	�C�3�qJ���L�1�y������Ѭ�G��m}!s��T~�wg�;4@&�~:�����7^4@�v�k�-���;=�'�hj���p�OF���3�p��k�Gzϰ��Ҽ�J��$lw�۬\�.��V��(��M��" ��2�����"�SY8��]xO�'��� E�7�����'���i���n)`�����M*�R-���ײk�dq4�	a<ڷ���Y���)�`וD �6&n�A�isހ�/F��p!�~���0�,�P(��A�ʄ��[B��Z!���~}L��	8P7DYЋnJ�:2鷤�e�6ͭh'�S^��6�kX�?����3�<f:��|ha��E�)�|�eK��A�<�$�#��) ��$�}s���`��O���\��E|�z=`VG=�J�Br�4Y�?L�A%������r�������q�p�%( �=��~�T6u�ˉ-~�%QB\R�)�7��F��,3Q�hTɫh�{1�= qŌ�F3���Pl�5�H%��R����ֆA�`W�ww�}����T���D���1�MF_�U�Dɷm +���n[�7LF�y3ŸY�Bm\*gC;�Lݠ�?v�aӪy�Ocx1*��G����f��M�~���.}��7 ޺]�$b<Pd����_����p������x��a�b������Bq%��f)�����|��r*d��ʋ[P�~)�D����tvj�ozә���O��f�����~�|�hm�w��-�O���IG3<�M��9
ju#Y��
5�KА��d$M=���P%�fG�,�'��?�/>��M�u��kӊ�$Zql�&XP��%�U�-῞��c�^�u����㶁^�xC��o7�yZ7�oKdG����ʴ�Z��o��mh�*����P{�J���0�s�^�̎�����\���S��)��ݕ<8i׾j��� �%��\�4�,����9&�:y���y(v%_�}\a���b�*V��%?��=��硛PrGHS��n�Z�/?p�4p����}n=�k���'[b����7+� �	t������t(g9N{��+R�� �!�!���L���r���D�V�sCN��->/�#*3�Ѣ�%�X
`Q#����$Kl��m�T�}!�IE�L��l�yV�=a��hTZ.�YS����A lT�Ru�4�g�*6�)���>�h׀
J��֕�C����h�r�V욊6qMŐy�VN>��L��!����a�xğ��|>$>`�h�/AZ�U!�73Z��|�GXc����;�=�5p�gd���۳-�����'C�t����NŵX�v�|oy	�q]�T=�?^ڙR3�����ݡ'�P�5��2 �oN�j&]DP(���#��iZ�fW�$M��RN&�'��R�X�`T�CX��ێ�Hqg%ހK�7D��o"�����}���:������e�$wa��M_V�>����z����t�������>`������e�Ng�;�h���zR1�$���3�9������F5B-�0��lL�2:��fZZ�9	؛������/�@�n+��}�oP���䓢LhԇS��A�Ҁ�:�'���^��R��c�ړ�c�#B�&�Aw�3��� i�߀a�����Hx��6�"�n$�sD�_���FVn�+�0�<�~�H���5F���Ӊe����I��l�,�郘��C�$!�v�[}�d@��I<����u���8�R�p&��e����_jL}M�&<��u�5�F�lL���r� �@���SE����_%k!�j2E� rI����ͽ<`�]5O���F n�W@�¤���dպ��ϒ.�Zъ@Z74���4���V?,?�<c��w�;��!%�&4Uc���RӋ`��pޫ�o&�V��q�ѭm����/&]��X��ȹ�:��z�կk�x߲�Kz�����cu<���U|��(�ΡJ��@��|�G��M�E�W����ȸ�c�.�SCS�U��C�x*W�!G���.�_?���Ʃ��wr7�����������^=��֌�9/�P��4.(/�I�D��jv5�2��'g�Z�x�p���w԰�?HSN��fXf�.�5N�L۪m�,�X�\�-t�c���]���A)����-
�M�$ѐkӅ���՞H?7a�|06��P}�dп�-
̉��a�]����$J����B�5@�k���[@ E='o�U�N3���4�i�7�8o�����v ��y��I�)��܎�.��*�G�q�<�����E�\K� ,���p����M��f�8�C�Ү��:xW�6��.�!f3��C�X�}���k%�O�O�"��|��#���#Q[�[��J��m�=��]�Z.�*�ŗ��S����]�l�[�p��.H��6�u�j���������g�c��=�|��1Mg��zs��5�t�"�B��WӼ(��H�����X�����a��h��[c�Xw���厦�9�l����m�o�T�ч��R��3�my�P�iA4��N׭��^�}6��5w''���ݦ��e��^��;�F��n��ׇ������.���\�փC��s�ec�\C��ժ;AЛןg�A8��t/N�0�ʎڴ����G�#�B!�`�}����a��m~�%���0bk�̕�B�x_���J��.�z޿�5����V�	p���E��7N��s���ט���g�@��=�}�NtRA�4��k%.p��۲cr#P�]"�������l#�<�hM����uJ�n���V�(�9#�`r<�Sg>��U�"JU�$�Rk��O�}4�sy|�(�ߌ�1&f��k�+'���mߥ-��w3�l����v(��#_	<�in�L_ x�Gr�ʄ˿Ce��iT�d���uGϼ�2�PQrݾi�7<Fp��s������_=ʣ�p��)�|[oy�����F':���%(����ԝy.�B�Lg�ΔA��V�6�!oG-\�L`��g=�I^!��2�,0o����=�u��~�(�2�swl���+�~��{���4"�^d�z�*Oh\�{�?#�4C�Vw��I[*<֯/����I�xS@DC�M�p�7��	�{�y=w�ǢC}gN���8�FaS��9C��Z�мh�H��7��p�	�y�H��qy�i�"TWV�P�ru��y%�NW9�'m�Cȏ��Є�i�X�p�Q�߃,<�d��>L	(�D�*_V�Z��#�K�>��Èr��k� �9��ċ@�V�U���ڄ��rݴ�:�BP��iF����(�4~n�c�q��Զ`a �tp��*R\�ov��/a�8}��4�\���a��Ҷ9��\q�s�w�p8����cBMtPՄd�d7o���c���4�r�� x�����pdv1�˚.�W�;@�@b54!d�s��`,�����\i�,�x��)��p4����c�'��(� wH
i�����p���F����z����i�>&I��qӨ;
�!�S[�Zpvcs�\r5��|�@�Z�]�M�մ�/EY���~�ldp*�%�&U}Ƅ��X���
�j�GΜ�^F%������!�N�w��`�[9ȟ��m��c�7�n��X�UP��P���9d�q�ޤu�i?��9P�S��ӪN� �ڰ�y�����B櫲��Ѳ�v�?��*2�e3��&ee�J�B-ŧ�<�U��>d~��w��+��	�,�10�.���{�^+�S��I��n��������S�덌V�V�~�� �3縮Vi��QX�!;4���z���;��[L����.��mp.��6��(Yy ����]�<�oe���u����i�,�DY��U^�_�]�vBļ�[����>=��Wu4�A^s`[{��:<��c�������F\.���(ks@�ؾ���q����w��cQ`R���Fn?+\�~���$�M�G�Row���Ӵ񪋽e$`��@���[��-�|1\!�"`�IWp|�4��D<R�� g6��Υ*�Y�����n�'�2��/�I��3g����g���^C�vY�t�}��}��y��)_�	'�����RcA:<]�ݲ  �.�3Q�f���A���M��K�x��j�����������Р���_[91)��f�֡��r1��6r���T��>aZ;�,P�le~n^���s���<.9��9�_��{���${���͘a%���D�(���� m���� �t�.Z�TK����/2��6�ٙ���9�r���ُ	��^PS���,�#)ҵf:��.�h��o�R�s�aϫ��M���S�=Z{7��ֳl�D�kZ��Y��m�?�w�Y���x���$��V��><��1��i�#%�8�mu�0��AI���ًg����%-�@��k�V6g��|.��c�����<���^��	���v�S��`�����|��YX�%��d���Fyg/N�V@���� ��_����zh/�#�صMlSk�J��"�h��遟�`������&8�U�d�GLJ�W���Zi�R�3f݃ }ET���Aה�.-�˴��%�=Ƚד��o�����oCi�S�"�����9���=�R����\T�aM�.���&� ���&��|�$[�^! �i���}��v>����/��:}���A �ȸ(Z�|�fnVM[��6�0)�Y/Ĺ6��S�9Zĥ�ص���?a��~�����p��`�b�e�%�azܗ?E���{ڈ�ej�+`B����x�xIO���p��.^�b>ޣ]X�����zC���x����2Z���'�/#a�V'�g��EH�r �uNc_�"^!��&TjE�~d��K]�|���SK�k'��9��Ep@3�.W�`�pV�#�3�q�j���N���^�:��\�D(�f|Њ� ��ޜM�`l0�4���Y6�T��a����O\t���*��@~�v�K��!�|�f�q0|=�`���B�Ր;&ƄaG	A&�h�@>f4��2u�����[_��!�����2*���*�i�3h?�V���M3�x��a���k�W55�G��́z��{��^�cY��ƭm�qy��fn����d��]��g��6�
Z�T�v#�H-`*�3�%t���Ρe��/m��fi r�lU������H=��E����HD��>��̾��NC�FAq��b�gx�<Y�o�1����/Y7�$�/ ���8�.�2t��w}��w5>-��̽a2͔,'v=܏k��{*BT68O7O�N����f��b�<X;�����׬�F�[���/��T�?R��a���`� ��"(�G����¸���U�x\�Y�.c��r����`Ն<���_�ߧ�1<L���k�`o��a�u\�D�r���0K�\m#x0&�P����������cF�/�C*Yg:*�����b^���B�9Nl�B'~�����(�֢��tn; ���(�lQHI`�&���dc�`h.Ӑ	l�A�c�y����3#&�XH�T�^U��K�0�t�e7��H��Z� %�^�O��|qs]r�>$5���,��o��B��I�"�4<�_���r N�7ނt��,3���U�>��񄴸�{����>!KcL��\e�M��@Q�]�)�^>�}.<u�׎�l�iw��+��_@@�!�W�����\�˚��"�S��aIj@\$?�'����aUث�! t��{�b����~F�䫡*;.=�hTU�^�Y#ѩ��d��9-��x	ҫ-���h�	{fU�n����D�.#��J���������	�SIFR�mcm�g[��&z�=U�h�h��
l"Ĵ+O��8�L�.�� �Y�'��X���&U[�:���+�Y�mʽ�#;���V���_�3�f��ܥT�b�w4�b��,��)޻j���E)��xޯ<�Y�`�%Y��d��ʨB$�T���]�4
�t�/ܔ) �l�O�7�qy����EN��0�ղ�~z�Uq���>Vn������O����n�I���?�8�W�)��8-,���.�U��\&� �o]*籾��>,z�#ȵڪ�;��u�/�R-m��&P�5p��P��������6o�s���"LeO�����~��������Knv��&�g��;������WOw�h�}���ʍ���
4fBA8j\�&��ܖi}��0k����!֗��"����$܊�L�6Ӧ=x����q#N�M%�"*�G���"M�"mx8�Yk���!(�3�|<(?�@X�.��zP-J�/Wz[yÞ��vú6N�ܳ ��x�������̸v�(�8ߦ�+�^j��X��\?#)Hj$.X�;:�]&��������e۫Uq��X�H�i�[2���(P�*��nv_R�^H�f�����>b��p�%d
�����Nڏ�����D��Ɂ,�_�v�ҕ����x�yG�k�z�S~���zc�Zr@s�l���\��!3�n���W�!�f�R����]�����N_m�	˨�m8~$87O�K7^?��cg{�3�
�[�j� �HM����i5���<��U4aZ���*�t��%#���9N���L��X�wtw(]�Nh�}T%SǺ��;��v�#+6���bI5�-e�(�v���/W�-B�A�m��%� J��eO��-*[��&�u][�B�'�J������ȿY}iV�ޛ,إ�晵��PLT
`s�����HV�m7}T�<皆�����`+�h�p�75��ɪ/��[����^�.���b�Z��_�R}�9b��F���V��Y��DjK��8;еN�Y ��h��(��Y�r ' �۪PS|H]����ey�n�n� �׃��N���;.RvO��kʣ�NS�i�yQ��/�cԴ#&UU��_7�:y�����Y�B��T��
��$��kv�n�
`w��7�=�|_�~Z'1D�M� �}�?"���rs
��;�HZ���Ћvu:g
��["�"uH��P`�a/=R/?7 ScQ3?�~͏�0��dd���	g�R-���tU,7Nyzʨy�?�������X:�\���)%��;�CE��X]=}��HFt��Z!��yU���0w��|6*jR�1����A����3���˗Nq�{7z�º��%B�'�>Kc4e���"F�b����+�vٷ̥�U�Vh�b�� T�Ĥ�zeBCIrNt��`�;�pM�/����R�����:H_�ś��o��|h��BU���#Q�/������0[���[��wr��ж̷�N	�����Mo�,b�؅�BF��#!l�W���_�0�~,�
;Lb}R�����?C#͵��án��B\P�����i�����:�B!��$\06A�l��hK`�ׂ�䳼�K�M&g��<�b���c�%u��N��������������c��>{�HW?�s؈�41�2�C�68���bg�q����G,t}vVP�����icn��?S,w�M^���'� ����]�0 ���ܔA��1�J>�3�<ҮY`U��:S��*
��5
V, �[�� �Wx�w<h��/s-�o�'(�c^7�?e�{�tR��}"��m�>��°/�#�;��S~�9o3��K	�LD!d"�׏F6����Œ�7�3���f�WPQ��C�3ݖ
N��'�g:�{gY�o���ղ�Z���K?���~�� �-q%��XAѦt�R\c��ii�G���|G���jY�
~�\��,AR��5�+J�y#�@����10��G䃂�<���9���aR���p�Ng�6�$��T�8��I�t�2��Xg��b��l:u��5:R?�� �Я��J�Z�s�=���'�H`;�jo�K\��L���pY=uz �Y	%�j���]�X �u��5��{6�pj���U��a'P%gk���E��%�T>:BR� �
����I�����U�����B�5o{kF��-F�n��;Z:�mp���-����N���>�)��kl��99;n�T|	z
���ߤ'Y�ۭeu���f]�����!����k
_9�*���#�cD��"�V�>]�i{�q��1��w	�||�7R7���� o�<�X���-��5�Ȓ��a��Sy���f���%)U*�+�Ŝ �u�0,��B��YE,��`6m׵v�v�J���bA�~9��U���[�Ͳ:ў����^og�-t?:
��,R'�`�O�Ď�t�hL��G� ����C���Re���0�n:
���K/�~T���Џ��5���k�W!/��o��l��#	jJ���N�#������
��#y���M�:)��H��WE�d�Di�f�2$ׇ�1�8��A&,��)<���tj*4$ŉm��9�un� �_�/�	�z{`���ٜ~W�.Vk���jC�zQ3����]�Rȩ`��)�F��/��{�ث$�kD�Vͱ��l,��S�/רn�w�����4������r���	b)�/�)�Jaz�����s�y��={�j��B/��O�Im슷���u���Q�ρ�9F��\c��Z�E��+()��>��a&ch���q;wa�I(lm�;���{�n#�X~��VX1�	��E��f���-B�a^�&�Ʉ�0��h���]|{�D�ڌ_��B��Ml4YXF���l��R�T�7��"�L/�G���n�2x�3N]l�5	J��nµ��ފ��@�Je'�xm����P%Z{��&Gӊ�ٯ���
O�=�P�o�.B���\t�*�>��h�hN"쾀�/��`��14�@B��ooX��ₙZ��(��㊷��Hk�1ʲ��\�lc����,��<�F{��JCւu'D�)����n5�<?:-�~�ج  L��Nb�㞄��3�S�P�#:�jt��ϑ�~[V�R�"����ub����������$<�]��!��O�;s�-����?��˷r@ց�JNr��yG������d��b���'��;��gFq�
G7M1�n?X? �z��xk�,��r�n&5��!���)$�X�{}���8�Ǐָ���	m����r%�>[����i�q�j2�X�g�Ê�&��Fɔ�{O��X@2��mn"!vָ,z�b��KQDT]mJGKu��jCE�^�6�_�K�n[9Л�8-����tS�\���Agm����X�0�0)k�;�-�]��i,��
V�K�#�t��Q�$�{pG�0b�z�0a�C~	��e%���dJڴ��uρ5��[0nW�F�4� `u����=���F�OIIY����dЋ�m讅�s�8�p�S�F�d��V��-��O3��b�PG�j�b�5������t�b0�$�
%v�@(�l����jc�}<X7y߈��?��P��E(�=W�$[����Дϸ�����SE����U&��B$������Q@�=T-{�K��_tH@�N�Q�_Vn�<�!��'���^!���٧~.a�ٗ�;�P��dFIs��`�-�M�D���� �~�o������uV��?wċY�O�u�_6�1�	5ｽI�m���
e�Ek^���l�-�z��rr��$j��BMA;�uJ� ��!���΂���j�T����
"��|n��QYÓ	[�v�0���&�{�C�k�j)�yE9�G��P;��D+����$�/H	�ɝ�'�&�M�Nu�8�ˣ��#���N��2"�N~^�&��6�t�4z�]+���	�������ܓ����Q��T�WC�o��"����1�s� '�Y"���
5�
~gtz�j=��~T�6P����P����XK���R�c�j��g[�����7�DA���J'D��rjŏZ/u���*�v�ۖ����oQ���T��N1^�D��s�X��0%^�Y9���_Kz�of�.y�b\�!�����Z����Bb�L�/���E>2��s�l�u8�Q=�2�_�/﫟��:0t��΍:��,N)�KrBS���)�Bp�Z�M ����]�X���J��Ҭ XZ�Xe*z�5w1���ew:��l�~rO>��Wv���f/e����RƚХm�Y5����N������߰ѕ
 �	�������/5#��"��0{�~�FD�mro��i�fSmOe�J��I���XY�:I�$�Y�Jm|��M���Y���:�$E���7��#ӱ�-Ż�M\�I��䧃(�� �Ӷ,�q��N*��tu�Ϙ� ���i��e�B�7��I�'X���(����-�(Cn�⧼ü�
,#��2���(2����-lĪ�y��j-�A^9Um��_�J�h;�Q�:�k�
��u��~u*�P�x{"ǃ�͆0��C���&��#�k�c]������ҋb�q��x�� ��7�P��!��h�Y�@���:�-qٖ,�S�L-
ᲬM�sX&�lm�|�5����w!^�1o�Ϩi՝�(%$�'�cK��|m�6Vޥ��q0K���I �p.��4���w���D��enY_4��-b���I����,u��͂�SG����Egz ȑT��o�l�����9'��d'qP���A`}��I#�/����&�~}>`�U���և�p�ߓ�uB%�0>:���aH��R�Z?\����e��@��?A��lk	�v��q�-]%�D�s5�l+�������?�(u5db�5t+�?H��F��D���U�wx�rL�g[ٗ���)�㹽��#��[݂�j��|�
!e's�d�F���& [!�ZO0��+&/�'�G"�[����SB�o�B���
W�zs���C�:\ߛ8�`�,3q6Tp��ݿ���4��m/�����݅�6���W��y�CQ�'�0@Π^ώ�ӿ*
B����{�A�.���
T�n\�an4?�j'|@������?ҏZ����ӥ�dk�O��X9�/3�UJ^?�/�5 ���݋��#F�1��+|���rLj$ńm.qz������~y1�j�EX�8i�)4D-�<a
��`w�B�M|d�A�"V��	�W*P<����qN�O�C*�/��1�W�0�J�<>*�T$��n��L<B�V@�-ʔ;�s.?�%�T�,1ђ*c:?{W��A�B�k����[��.Y�g �xC�� �6RJ
6a�B�m6�3���|���h��dΞ��NA��Oo�u��$z{>��R(�D ���3�rD�\�4F{,��IZ#ﮑq@����W*ܚ���шӟti�F��D�d��׏4��0� _�U���M�H�2����;M�ce���.���wQ\�|x�,�����4�dj䬓��Mx ����j}�CSk��L�xtj?d oܹ���Zl��`���O�]�Lй�v��W��
ג�}y�o)lSu�0��<%���}#`�B��h��#���+��Xv���pdJ��֘�sLTyD�|��ԡ�W~Ô�I��H&� ǥ^��Ӧ˭�{�SV�
��������o��o�^�04��1!���Ml�4����;�#}��dDmXo�����/��N#�h�䵽���\y�6���6�II�N4�.'L��c�G6��<0[���i�e�\vl����{7��E|���5�`[�|�u;'N��t��z�t1�i���~`���$<{��hݮ�Lpl����5�Oy8E׬�@1o�{A%��^��Lq���8t�l[�N
�������hDȨK����b�m��N"���ͤ}K<z�,~��ݟ��T�_�^j�BZ�(��}4K"��_���M}ڨ���?��Oz��m�k0\j�<&�lX?�9ZT��=xڦ$�0�FW�S,�}�0�Zc6���{t��:`5��0��r��z:��_�W�t��D'�BeDn�?�"k��+X�4�w#�@V&G�#���@s<h��vBe PYQ p/��>L���Vʃ�+H�)_�b��h���XsW?�dp:��TJ������8��,�@f Z����:���h?� 5��A��/2���i�Ž�M�`�#���K�OVg���2��h���ύ�ң ���~j�b(]o�VZ`���{x����c%?gD;vw���;�%c�t�3U����7=��P�v�T��h�&F��o���~oDn�}h�"xT� t����/c�M>T��Cpl�ڪ
x!T��=�f�G}�X Z!�ƭ�I�7�O�ɏz7����o���E��(���J�="T;�Pc�`�(F�g�88��3���L��(B�^��VN)<D�ʯ�f,Vb���R�!�:� HF�7�lG�9o��Eu�F��w"��@)�>������;����a�w�#�+�w4�ƋG�Ӄ�蘷�գ�5>����@�M-.h�:�Is�M~���$���ۛ�4��:�����B況ǂE�ϫes3��׮ ��Vے��Gg#�nD��Y�"��g�n�v�� Z	"��¬Ꙙ�O��m�5��]������M1'�욝�a(�YXжhRB�Mm�<��KY9�1o,Y�U�n�OeI��XK��Ŏ����\~�^�&�V�	�6uy{�R]l�x�r1����?i9!@��{MXr���>th�?��EzW��O��4�VK �\�B�uU���6� d�3sW�OV��.�+���>l)rH���j�Ͻ�:q;�ql�եc,�f��[Һ;\֦�1����N���l�;�6�N?+c����W���#^�C1��,��Q��GI/�Z�Xgr�p����0����(�AV�қo�N�|�ӦG�]��@�˧�fT���em�ԄX��lZ��-�b��l<o��笶��� 졦�t�p�| �JÊ������y�B�XȒ�r�`����jX?V��N։����]@� _1#h�{c�X �?`k0-N��]
	䶬$uhB�:\:�!Kl��EܻlV��:�,��7���W�Ƥa#��64���.�Tɲg�<b��4����TN�ήc%�a�H=^�����Sh���	�̋ڒ��("z�IN8	�a ��)�EC̋MV
	w�ŭ��"ŰY�*�XJo���ڽ<Iߜe���a�%*d����pӆ���A�zf����1{C�ЅX����O�xn�FX�ܚ����B�g\d�Y��0K�yj�?��F���+)�1$��ڃF��-BЧ��(\�Ex��}���k�8�Z��-r�s~
��5x�У�Q�~���S�{��(�!�)�qx-q�f5�VQ��4�炦����&ˍV��g�PR`����	xFQ*�>{w���63�T���ͺэ���������"�C��_�?p0��R���3T���KNw���(L�Pd�^�H
��"�.�=�6�|�� &�hZ���q噗�t��g ����{'�c�#\=���8�G�Ͱk��7���mx�U�}��^HWS]ƏK���!��G�M.E.�Y��&�E��k�֝�E8��N�'���K�t��Â�Ͳ���ޠ�l���m+�Ul���|�]6\h4*2+H��|�U�W�t���d� ��D|�'ǹ\w�J��E5�r@xY���,^j=#�'��t3q���1'��T�(-�8��p���X�^���.#{;�劥���j���OՋw��LW}�-�a��t����!�Q6ۙ����;��*וm\���&Q�vS�8骿�T��	;��s L	�O�`�l.�KH�I��5,�Ϛ9���\�;u�^IT���֑�qA��%jD>����Sm�\ �#��$����F8��xpu�RS�q� =�b�9�� HwV��78jE'�1��#2i�����Qu�iL�9�_�ۄ�L�ή�PC�|�:0SC��r�xr�关t*p`"�����68GZMO��%�����P�«�ۃ�F��~�G���K�|�~��`�ꉛ�)����TY�{oUo��b�49$p�5�:-����5`sN���c���;6�$X�������_�������@Y�m����f@T>�հ��yF�-����r$*U�0�@
��w5�g{,��Z:Ԑ���zv#��
�s3;3�V�~�
<�%( {�h�����n�����.eƸ-�Xla� �D��FZ�R�������)��M�2 9;a�t�dȑ�of��&��S��k=����U ���m������lΡ�\�17��$��M����N��
�z]���{0,}ϑy�G��jҳ]���Jhm&F^�Ye�$l��\�M���e��%=G89����s��="�HP���3��T��襌[�+�W�>)oOebfk��I�Y�ŧ��+�Ő-����/�$���ޖ���a���E	,E���ǚ��4]�#�v>�0�Bpz�VG(@h��1�B��W�@]]�G������7���N`����'��D�	)�����mה>��U������,�Дǖ�b���.!�N>��Q��0.��7�(����t����@R^�e�zV�^�c�����c{�'��r/Um
���4��L)C�6����"�[���5g�C��j���5STOh<����U|n�P���D��Pza�p����[ (B-폈�?S����}�}��N��F�L�F&��U����� 3�r���SR���[[���g]RY6�:�7)�$L�F�&#� -�EOneO�����	i-�\!�	��)-|���@�=���^���"�_,�15e��0���	TF\z��'};�9�����tG.d�Gc� ���k��4Ϩ(�*?���Җ#0kWY�}|UY��c�lة�z|S���7g[����:|R�f{����Hm)%�D��P�
Q2�".��8��]c�:]�>[�y$��5�$��B�IG[�I��C��̯���������(��d�j/'�f��k�E�u8�ϛ�X�XYY�.�q��������;t!�,�ukT*�m���B��qhM�/u5,t��!��C;�VJ�s�3!��l���HA��40�L�^�%�. �Tԯ�_��iv_M.B��-򋬘����mGau# 0��;|k�%�[�+óki7D��� �� z��7uAc�&��:�~�3�'��#�����
�X����_i�X�ܠ�n5��A�ckN��Iӊ�ђ�8h�
o9�x�������n��n�C�M����·�W)
��:�)o��_���z�O�l���+�iV��0��l�B�d�V7��P��$:���$��X��Li,�����r���@��t��U�(�M�=>`$?�6.A%���N���>!�ac��	Y� y�Ҩ�ʑhk�bL�?�0����o=̠Z���@���L����3����;Q����d�.��
��~%7Ċ]�ԙ����Z;���U��7����:_x��)w��w����������{-/υ)�(i�E�C�8Y�jo4J�U�d�g9�q?����W+�Q���J�39ёÓR���x��`�6�C���>��('�C Bo��&6�9.��_+'j8Ţ�n~`W�t~��e0�.1@�	�p��uo����יt�#ml����ov��sYy��W<7�Q�ǯ#y?u�Y�g�L:��S�=寧�p�;�OR@�
���v��NÈ�g��.�^���]=uo7W������P&�
��:��覻CM��"�/	TJ�w��K���8� ����"()��o�|{����n΃έ_�g`p׻:�'���������?mT�j��[�M^x��_$|~��#�f T�>�k	��-hM���Gw�t�@�G�+|:W��%=f��Z����4��?���фigɱ�N>�vZ0Z��?��:x=7b%	�	���%�����L���R��-U{����A�e�����e�`V�.�Z�M��U&�g��x�P4^(�8��7�Z���E3�<ur��v�b�(�mK�ϣOa�H��=H��T�,�S-��7EBc��v�V%MH���GC��7ðے��n�r�FLA&8s�'ĳ���T���Ŕ��)͚��Q���B�r��F���A���gpZ���pES
CG�b�oh�f�Uʺ�j��EZB��Lm��
)F��fq�k�X���6����NJn����x>�ao':$�(#(�'Ư��|�j�X�Y�]�k�|:��)'O���Ng�M�YQ�y��ę��\�6$c��o$n��.&�d��a�r؉�,d/]�jU;-��5}s�A=�Op�@WvE��*y~T�6K��'[6�M�pwPh�r���0z��<�L�����c)]�p�����{�w{]\^�[��h�na��~�NKi���K��TBmyb�rgѧ0uO��['e�!���8�����%i���j�t=;�й��U�������Jbgao�ڵ�9�U�V��=Z.��{��Y��c�h���R�O�-N8�i��U	��5�5�n�Ҷ���(l���!,�yQ)�*@e^���y�?���d �:������ꟸ���Ҍ�FXO^ޓ�O��3W6�U#�l�Xu�qn�pL��R�������x#N;�]� y�,wLE
 5�ܽ���)�[�j�(+�h7u*����[�*�h���3?���_ķ�cl��PZy��e�ٴX��JZ�Ί]U?$p@;�/[�M�J�A�2�RZ������� X����
$qs���\���($�Ɛz;O�r���m]�vτo��掊�{+���íV"Č�q�'{�l���z�r���g��͖2���b��w���vQMØ�Bo'���@x]�qx������۶��W��O���,1��ۥ�K�46Lo;�dB����2<��06�}|A,�B���������$��*yǗ����`f�0���=ۅ�N����E�G���G�&^�2��	O~������qў���n=�L��_;�S�D��FU��a�J�yD`:�A���N��Ǵf2(h~R&@��%���	d�H��[gq��Y ��׊�������Vf�">\[����tjl�H�_��i��=�(8Z|���ò�*��c����w��X(߅J��w���9Oޤ��΁����C�/��(��K$SsPS4��rH���6g͉��o���)�P��/���|����]�-�IW�D_��d�>���I�C�鳤n6���A�S�r'` H��/�`�e�?Rʑ���|ٞZ��x�Te���vِ�b�I����i��U�N���n4s�2�D���iŪӆ�$0rG9.vJ�h�~�9<p�M�����!!뺡YQ\��>��Q(�H0�/j��Hz�jf��BD��͵xP)���~�*a����S$Wsy��F�c��:���>�|�ϒ����g�˞��<,A��<#I+���{����w�A�Nw��~�^�g��� �(�M,�aVE'.��@�����&pq�b���H@q����Az�=�ԧ���&�V+�V`��,?sJ0��낯�Yم=ͤ�N�bt+[���J�!L�)�‹��x��q�T�wkRjH�߁EWd�� :L�k�Ɩ���$���������3�o}��/e��� ����B���I�P�R��F4.ͦ���c��a��$dd�	�PrXr��ձ�D�5���Dɗ�?��>)5�;ޮ:�>����D�೰x�E�ĭ� ��x������QЏ�-�F!Ce׵�{9��eof-W �B2�2�� ����"f����h���L�`@�؁@�6B�!Ю�ڭ>�Et�]�ɂ���V�ŊT�d����\�dE6U��Ȉ�q���D��gfO������R�,�S�ٚBTXnlľ���aӓ�;Lw:^��^J_kБ�N�3ۓP�v�� (5З,k{aс�֧��.}��"-���O���e���\=����X\I{����S������M��Û���宰��ը���JIW�nИ.�	cĽ�e�������]X{�/1?��R�h:Ӌ�fVT�:��!�����?=X"EĸL�Fp*?�[����2�;٧�L�.���ջ�����z�>���W��>,fd�g�����ud6�R�ͽ:�?���z���{�2ИK��x2!��6� 579��۰	���`�����;�v+#�6� ���"�1e��=I)��(������u�n��*K�X[�;_A�<��n���b�i_��P��M<��m;�{��]\E�Χ�c��#`N _�x�e�sH��sc	��4ԭ�1��t����<|HM�I]!�,�s�y=~�7NS�;:d=���k`�s���qzɲgx��n�����!�G�ʺŖPv�EH��~"4���Bu�T��t���[��?�
�o&f�Wc��[�-/\yۅ"
"9����c�t��v��*W?F`�ű�ySXv5�� ��n?�T�]����1�gq�D'�H{�l!U�E�.w��qp�5�`��<q��O����5���A��UGJঢ়����v��w��oX���yG�6�2;O��F�������wF�T}��귺�*�N�� � ���������ΐ��BΊ�Fi�e����R~�����cG��l�\a�9�t�߬c%U�F94�YR���2?<n��V'����ykL;o�]���&�-�	�`�\�ڔ%SⱭ�И�T��{Y�i�%�0�OТ�Ec��,�ɀ�s�e�i��&��co�s)y`��SF_(����;f��C77?��y��j�l�f3? ��dJ�GW־�K�ׇw��GUY���;��չ���:�>^��ї*��2�"S���@�d �� �hF�V���ڔ���ŕ�Ǭ�&��]Ӫᮧ+����9F��pg~ϟr��SkwI�G ���Q��o��bq��SHlK��k㦉�ܾ���}�i^_F��k��ki�����Y~Xt��H�k0�R&ю�~���4J׍��":��� �*����id�l�c?���V>��>1K"�+d����=�޲:Z�hx}CE_��d�wB�n��`|s�9��w��U�1J��76���+O�+'��lِs�c��Md�z�e�ˡ"����tC�V�T���y����X����� ��,�Z�r�^]�vG���O���m3m�5�����@��ƀ��Oz�����F!���]����c��{��={��k�v���O��r�y�ڞ�����3�l�P�,���Q���+ݸ�x��=�vXx��o�����\DL�pamm�%g��9M�ۍ��~�6f��(2��r��-^"��p妦�K��1�Ⱥb<dM$� *<1��H0���GnA�a�����o/�꺉���:�\���������I�<��Z'F*�r\?����O��p�=t���08��͜�03��y!k_Fwۚkw���ԑ�³�8����[1�`9ܾǂ�éAϙ����tz�����-���z���AړA"b��T|8��29�LH���EJN��)�j���.++�=4y��������w�m��\��?���@�b��b)�,�u?hT�w"</?��Ӟ-�����Y�زR�#��/�v,���������P�O��&Q���]^�)"��u�@d3�/"�GI�=���E:�����ds���,F1c����xـ��cQ��+�lz06@*+�O��N��&�i�˼xS��RG��n��bxC7�=7f�?�eػw*6����en8:G䣌M�ӏ�hQ_�B�Of����o��+P�����Miɤuv��7�~��3Y0h�A��oꢒ�T���W��6�����h[_�� mi�Ç�M��=�1� � K;���+.�[NS�����t
^�H�C�tW���d�:�G�`��g:��s*��q�?H�p6���@����%j���Z��m4,�rp�6Q�H�7�g��Ǎ�ߴ���d���8b�"��J�.�y(�qɸ�Q�Nj˕�mH3�k�.�m�0���&|0Tl�LJ�6��z>��MR��*�����p��E���Wxj7�e���g��<���Hg0���
A�ԍM��b�ʠ���{q?�0n>Љ0��,�o��$,cyMa��Ẃh���6:���2}���!��$<Qx�{#���KZ��g��ɇ<�A>�q����{����SE��չ>szD���2�!>�J��Ȑ��$�2#x�&���͡.Ma"癫� hi��6�^$`�np'��-J������O�N�N��C��cc��&�D
[3���ǤB)e�N�zBjqH�ū9�� �J}) �;̧)�j?��#���#���ŏB� �q�����k������qV���+����ZN����!�;gʇL��>!�`;�FaՕ^"��\O9�@�L�ٞ�}O��O�[�����Y�9h�i��ԕ����d\��j%Zu�ݗ9OwK���-�C$[�(��7ˆ�tV���~C��Ocݴ���:�N�Y�k�)(����><����0^��%��*�[%��k̀Z�mT��J��5�P)
7�-�X��tҶ�YU]��>�5W��| ��7��k���@��G����ل¡�0#��({���5̎�<ڀBl�|��M�#�5��<��~w��U��By`I�:�͌�oJE-!�`���z��f���qyj�"8���<�zIac-Ve`�o��-��'1DMze7x�'yQO���B�mG�?�_h`�x����6�Ϻ���4w������?�{h�s�M)F|�v�.=Bk1Qj�Ge�_�R�[`ZNtm��
���H)����mh�#�k��,�0���!s #�ȃ�;�'�Z���a��[
��)ڎ��N������1&��!�%Hb��T���m�:�U���G�9?/�ir��x�S�n�c�;l&%���Dɍ�l���v-�w�Q �ė<���Z�Y����p��2���o������P�A�G���x����U!.�L�z��zA�LL3�|���N/QҮ���Dǖ��&v�K�׆�y �K�([B�Q-���p�Z�]���LY�� �o�-�G��Q?�9���GőJ�NR&]���X��=�U��b��,a�F��`ї��/�p��;�����f���7o��(�)a��(��]���_r�q���9*]��i|��O�������صH V��I0�O����g'/S����YH�EX�+�T��;X�5#��ū�޹�Y�r6sf�mS$�����X@���ǔ�~1yF����^�K)�e> DE�T���������.Q>aG�}���,mG��RCpK�'�˔O��ν��e���S�(�����n�QH���o ��a��R��3Wp�ܕ)��gB�ζ��~=��u���z��Z�>�U�$`�T��W��.����\3����"7ɴ����)v��F�1j%�g)Ih�jw�����`
D1��%KI-�)Nq��N��$}H�������=t�*�#L�_H�i���bDa��%^f��1C]�����U|�l-�PÄ���*��jl޺�>��d�w2T��ЋK�_�R����r�.cNi�b`oi]UGf�k3��,���,�T�#�X�E�&�&j������u��M
��*�<��s��׻䍜#�hQ ����1+©-nf[�Ւ�u�\�+�5�R���
󇹧������'٬�oo�,��TVp�>�{���M�����w�v�fO���;GT�Z��bc��=CgY�x�ql�G�B)`DF��i>����Lj��ێ��&��gw����.��r'���Ϸ���������ҋ�z��ATV+Fq+�S�����1O���v�m_���\	Jq��Kg������=x)M���Bv(�LO�)[�\���rLu�w~t�؀�N��)�c�=�6�d�C��1i��&�����P��8���'�S4FV�V����1�S� o�8�g���E�d�F.���׈� ���x�Dg�\���S�da�����1�s��^ۑ�4~��]�J��q�gC��J5�{x�h�a�aⷯ�����N�����QWK�sH苎E���@|�$�`���pWn��1ʏ��ۜd�'ݽs<�!��[�Q���j{���M��˛�"�`�m����Mr�B��T:5ӥ����Nj��\I�Ɩd�A���X�X�4��F���h�	�F
���-�Bf�b!"P��f��S?"@��8T����O�|<xΠ�M������/W�qS3�{<����H�a�_k����'���־�q��k\s��f �x�;g����~ۖ�a�j�7�d��"��JD���;�k��Fgdl�P�jE5�4��Mn�Ŀ��V�������@�+��E�.���1�[������X�nܕR�H����zh��Bb�׃��O_m��W$d����=����"(�MJ���K=wvӻ�id��NJB���^�{$�N��g�K�zT��9x�&z��	�b�y��JL�x����6��S��P�K�b>����ڔ����B ����<�H������(�
�>s�����y> Hk������4�<t��
�ppĬQa�A�s�3k�#��@�<�����,�+z&���9�+��)+�A����%XX��Yy�Z�_��P�&L%���pނ�{�67}xQe�6Q�wVƨ����j\�'5�mYO��}o����ڨv?���7��t��z�ʧ����߭2~;����Rx�-�o�~R��g�o�J8w�Tn�I�o�:Z�K�_"6��[�p��?@o������HA�RV͘��_�M�!�c�c� �Aj+��
	Vw�x!o3�Q��'��<4`��i\J�w��`�\�{~�u��N�$�ed�0��NA�F���z]|Z2�1:	��,4Ҫ�w���c��ܕ.�q3��/�i
�Q9-=7~����i�V�I^q�}3����ߣ<�)��o���F�G�1��m�d�=�C�wP9&ȡ\k�¤bY�som���x����n����t�)�mB���z�
����R<���F=<Hje�\k��>_3��i�dS�ƟG������p�br��/�콎i�B���dk�t�%�ژ��0ó���ս�F���/Kq��bń����R;[�����Cz9�nMb����z]�Q�Qү����E�7����Fܿ�5�b�m�	������ݣ���B�(�~#죀WD�
1���ձ���>�nINn�p��m�ހ���%l��b�ߴ���L(���_T�mx�t�?w�w1aR5�̚8�XUW/j��-%^���_�f���9�)	j�hB�W�a�/��4�g���lӍ�$��o��x���GvPD0���M�E�R�Dol�@njs��N�Z�=j?�=��L���鈟 -o �)g$�_a+�5�����s@,(zNc7�U�A��a�ޜ�懼�32�8R;!�������M*!�{�R���,���Q����1q�	󯚙��.���?�����  A��|�ɸ��7a.b�B��֗�BuV�9��f��i'��,��^��%B��Ye31yѶɵ�ƪ�N��n��V� є����o�65��N%`pb��Rb���}+�#s������zpGC[�3���XC��|��y�b�j�ξ�`�ɤ�����q�`�{�Y
6K��"����@�{���R���{�)��.��M-�)�v�H*�n.�TD7��b�i�hO�o��Lg���>Z�!���õ}�PW�9*i[Ȅ�ƎK�H�fj�����yx��!sI~^nr/��i��l����	L4i��a+�c;V���Ƞ6c�^
h�M���ᭇ���)��׼�-:˭,nK`dR�x\�{aE�-"P�]+�6j36� ���8Q�ǰ��4)�Kg;��b=�U2� ܝB>�W�෺��`!C�eA ��?r{�������>��f:�?��
vH�����Wr++�N4P�wr#u �����,>�8��x�d�G�����)�_��)� ��V�<:��J8�dڱJ�0ҷ���Tjy %��L�����ٝ�>7�������+9�d��ʏ�O�2�� �D*���B�	��̶ߒ��{@�LҌ��yf)��??���<?a�짬�}�N�8����[�����)P��z%���G�K�q�cM#���xX
�c�Gz���3�wR,�Mb�Rn��)���'�m��h��w@옒����)3��q�8��������}.v` �<ؘ�o4�r��������j�k:E#J���%���Q!@���"ҁ�(�6Ԩ�ӄ8g���j���L3	�Q+Eoo��A�%��V�m���ꇺ��������sJ�п��L��ak�!F;��,6��̍��Dg�I}����~'8�&���|��}�����=Q�+�����(��J�!TވEQ�ewJ�y��Y��������H?ja��0C�}�R�~�->Ʊ�By�'qG�e� �����f��J�A�rA���}�/�S�&*I�f�u��R�gE+�D{�BN�S_JFݜ ~6�(@E��E�5O�-�ѿo�ҡ��l���\n�}�W������-#���q����_�e�B?&m�tmWj�3!�'�@j%��fv�m���B|�AM�ֻP�J�vjHǟ����H�A�9�Ce=��*g����>m����R�+`n,�g�i[ފRB��-W��_��1Bm��(���?]{G�H����T8��z-��ަ7iMa
��˫]�n��t�!;��ſ����#�+K���2�n/�L��v����?��O���G���9�WL��C�����ʥ��)��^�p9f�ϧ�g���N���bH �Z�+w�:�Ȱ\x���`w����+�	�y3]��xH6������iK��ԶT6�^�S��p�dc���-_���=���c�t�^c�s�\��װ�����%�$�	��j�J��U��u|k(�O��NG}�G�Y�ںtǱs��9�ц����3ў��0���Oe�M�?���:	Mi4�)]�eM2i��k,�a[L|ݷ/YW��oh�Z1��&�y���va�>���/�c*�MDVq�����w�xv�9n�e���YC���������k��$�����@f�8��xQ����y�J]�F���ZЅ���G&0�p��*%d�L��}���4vxs��3��?��e�i����i�Лq���;ۋ4#�N��Q�5mj�t���RbΔE��{��t����J�1�1����g��$�����ʍ�k�ހ�e��W����?���! ��7�N:j���/]
��=y._̨իF�� 5�����퇲��eC�Y��[Ji>��x!po�����rmr�A7�����W��OA$� :���d�F`t1fJ��5 {��T�t��O^���ڡ���>C"��n�S&�G���^޴�Q��W�Uj�G+Z��O@ z�@�o��R�^JPx��2��h���LsUKX�+`�y �"�H?Jt�H���q�ߢV�<l�O���H6��9$�G;5�_��2}A���iX(���i
^*vq)6KF�B+'���Xqa�눦}��E�WBx�pjG��L����r�Ο2hT��*g�q u'�Gt�;��
E�R�2���t9�;[{Qk��Η"�g)� N��)����g;4&Q,�� e HoWQ8�v��7�y�%#?��yWf��w��*�~- �Ӛ�V�F���qr�ω�ں2��	7t�^��aD@˥9���%���s�������Cy��߽M��eA�$X�v
wQ+B���2K� �b���ЎG��Z��^�|p)�#l�m��-�[�
�,f�s��J�5��7��\�V�A9����PvIE4X�D���qȞs�D�ȈdN��P:�o�b�g�_�DV��~$�D��&��)��U�W�~/�A�� f���:8���P�͝nDPb,��������p0&�cV���&r�Ҫ$"���#����u�?��y�k�
��Y�F�)9����HAY;Ap|'�dS�.���?�ܷ���n

�����.S�5f���@Y����#
����>� +� �v+�yR�E��i�b}��	��7⼵�0R��fS�:��Y�[�����	zs��gN�3�_κ����{�����i9�4Q�[��u���ӽ��0_�H�*�|$�56nT�CD��>��E*�M��'J��Kg
�YQ�Z>�+2)N
Z*Ike*�l5_���î�=)�M.�y� #PtԎ�@�n���,�
-���{S�T��+4�J`	��Pk���b�$�?r�\��K���A0K/3��~�w9	X[{rZ`�#�5W�;-f����xѰc�x6t4��_���7x+y�����w�2viw�:�h�:����N[4>S1�țϔ�d�]4fh�X�KI�P!"ض���o���
�Ɂ"yR��b�L����hl����}��ǩh��b��n�@��׮:���	���qGU��%�Z��5V�0�(^�	�6��!�[e�������.pO�f�J�k�@N��i�s��E�Ӛ������IE�������/	�	XC����|Z0������	�T�O�� 0P�w��璞�ܸWt*�l0`���m{��m��_�I����XV^o��7���oQnp�UAR?V�����pORE�a{B��sC����J}�a�:�L�#�Yӫ�@mp�W'�����ăǗ�me�ω���~~�N�p+	S,O��7Q�dn������p����Z��{"{���lP^��G	L�������u I����G��_��Y*Q��;� ��O�����ᕆ��ʊ�^���S�l,Kp��E��R��2����Ű�e�ץ��,��a�����%�*_m�k�q8��G�ޜ�D?L�A0z�Ll�������eB'N�L`ڠ 5t~�zW�_K�qQ	
$o�a�0 H�s��v��?Qs���JЊ<�}�{�dbO�R�v�P6V��7�>e�H�'��+m�-����̬P���r�a�� �"�~�5��P�[Oy�в�&�4d ��ib�"�d�F|sJ�|41W��t+��;����!�h˜%.�]>w.g3/\�Ġ�#)��i[�KKS 5|�A������C+z*Nڻ��J�UO��I�����z���[��,��2��7皣�_�t�R�����;szZW���p���a%�k�V����d>T:��VT���v�B}X���v�N���m��Ic�ÅP�K'Ty��*�R.���g��Y���*g�"U|�N� ����w�^.f�56fp���踇��ؗp>/e����eA]�ׁ)\u��1��^�$*:]����_�6��X�u�u�/�o�2֥q�]j�yh�D�Z��4�kڽ�ϯ��Q��͎��{6&�#��+��X����{X�m�i�7Z�j &��Fm����Ǳ�Ո!E[�a
"sZ���?zrH�f��iF��C%��2���v�c��.�>ϛ��e��o˦�<{_}�?�c���o�S	o��!Q8��W�~K�iq��:s�z^N'��#����bRy�Ⱥ��ͼ��K�'��{��2?�Jrx!��䎛�sk��³������ѿH�{�뤌�n%��3�e��N�N�T�T5���UH�#�����K�,�36���7��3-~���鳿Q���p�,ReK���4?�C�Y�.���V�\C�?"'݄V�WD�k��L�{��@�]�F�$ZZQrp��*/�RB3 �o�~�{}|Z~m������Jc,{-�1%�I��+�H8�11�h�:�o���;��\',�ϟ�N�!�S4������e���S�q�w,�i�QC��['�.G�j(�gF?R�ߒ׃��~ݰ�2��q˰���^t��پK����O�ס§���a��2���?�᭶ƽV)�����h_Q ����}�Ng�3�Q�DޚF�}??N��#;���U��a8B~e�e�M��ܿ�+�c��s��y�V�-���ب\�		��yu-�Y���0x��g��e�d��׾̈6X���C�W��>��nW���qm*F�f!N�lԯ$ ���7h�\�I�<��[9m0��ߌ}������)4u~��.����7�ɤ`�4�·b��0�H�[?���O���4�s��:�v�I�R���ARS���#s�]�ѐ1��UZ(?x��P�>_�(	s��O7H��G�<�'o_D��*���������UC�\g�c����-��oٯR<N�$d�!��G���%�P�bÓ�yi*cu��� u�͝�iؚV2x�~�xPc)�z4�Y��qq��y�Z''��"}}���~�M�o�U�v E�H0�0eQ�N6�j|Q��$��^����/^a�Η�Vf�t��t{����B����Z(�9�9�]�����+ cS�AqF���8�6��Q�N��B������XI�)�D�J�-��L�0ߍ�8(���M�:���h�)�׌���ur-a����vZ�B⎕D���瘠a=A�&�E0���4�ƛ�[�5 �{��� ��,g�;Ϧ�1�Ǒ����~c	��8b�&��m���Oll��$3��lN�fU8�Q���z^ʐ�g������&;-��t������倶�A����f���?�p�i|�����7��+����~��f*W��a�@���4��1]���Uh���d��%k�6W�uPZ�v�з̠_b�+��A�!��3�0ny�K�X�3{.�Q�khDú������� �Rz2Ƨs�/�VPH �,/��%9v�3ɢ��M�&�j�FV���Q&�`4���W�ܰC�"���ꄅ�%�0���1��Dk���4��m�4��LQ�&z+����՘���^o��]H�D;�����J�o�Mh`��þ9Y"�@�s8�!���#�	��N0k�g�^g��`Y����>�|r�J��l���b��SO�iC����I�ޘ{"��GM�͛���� �t��N�cSO\��$΍HpR��OJRw��d�<�z|�Q�Z
���f������N���;���}��3|	����O�xiֵY,*��u�naB`3�'�֊;	w{ue�*��t��	��"�qQ�d�1E�װ�O�a�Ld�yBKUm�^�F0B�idCZ��icE��h�"Ŏ��]@�)�g'������R��XI�F�n*�<{1â��CX���!$ `�t�#��JFC���c������# �F�x�7pĒ�ߒ{��֑%�|PJ	�/~G�3}g���X=Ot�-&qǱ��{?�M4��!a�~is�RK�� �»�=�����Q�J)N#tnb;���oF�Qe��>�L}�Ꝺ^����?�%x��A�����K�+������	y{��H@��3��gņȃ�c�8�f�M�8����m�R:E�@�Z�����!U1ć4D+iW��bǱ"t����m����_��.�Jܾ/`6�Q�K��G ���a:��p���l�pV��;�ϫ3�+�,�v�O�?�z�C[%��x喋Aڟ�ߦ9��o7@3�����b|>���7n��q�2��j���6�C7T%P����m���q�V`�u�^B�lY���Y _�F���
�̑�c���|$7=�́���P� �<&��/<�������_s�:r4-Yj�5�E
O�;e5����@��e͞L�v�`	ȹ3��-�t,�~�`�Gȋ
�{��,�x�oW0����+p��7�h�4��e���]R���J�?�	c�^�/��.�b����H9M����浙r�I�
i$͐��NÏt�C��<N��կ�(�&����*�5�?�]�m�:\��xU�x�{PWX7��+��׌=�i�%��e�4{��W��oj&@�Ε�-��1#Y��7�I")���2�+qx.nx<| �:�R�/���8´��$dw���eSP7�c�L��"�H��bq�y�0/%��V��敧7 u#���H���"1C��9�l^��ӫ�u\�_"�ߓ��ؗ!�8j(*�^Tu�!�W��#�Z#�աɺ�^��T���(&�R	I�N:qp��ij���r�L�1����LR��+�eq)�E��?"$(MwG��#)D���G� ��<�/�Q1f�a?�v��TQ�U�O"e��ґ��t��mp����#���҅� �X����x
`�7%�޾��+��廟$zt�l���"͞����J�_�f��7��(�����z���rƌ���$��l%�u}ej6�?8��d�	P6�'N>[U�/K= &��m4b�������f����Yy%��V|n��0�	:�p��#����ł+W^�'X�Y��h��r�c��<�5�Į\N��"ʻN6�j���Q9�Q���¤��iĞ���d��sD����*譫����B�W�n���TF8}�~���5�M�K6N�yJ�>�:��x���5�´C���Ӥ���43�����n�͖E����b����Ay��)UeŒĝ${l����'Uժ����FG��ç��!]ށ/��;�����D����<Z���d�B�xFO��*��^�.掂�:��DM|��C,�1kq��z���	�;�p�Q����&�����r'uO'�Έ<�Rv����o&� ���PSމ8<5��W%�of�=�(�e�e��L���7��H͢"Q�B�ܵ�]��Չg<<�����ik"3������A.$.�H.�1���f�  �x)�]�@_x�l���
�k#��{0�`����X	]�����:�3��_׽�ڥ���b�LֵdN��H֗{:B��8����HLc���6�*�J\�.��W`l�r1;���8bI��Op+�����^�Ë�0%,+f|�ѿw*S��j�.��c�"*�|�2"��[i�FK�8J�[*/T1���	���$)�ƨz�g_@|�%�m��ֽc��g�_`�s���`f�i�jM|�n_�\��'Wĉ�C�Տ��dl��!�a���ޖj�?��Mv=��OY��5�	�dv1�˜�S˰�*:�O֨�O`��)�L ����@��Eǁ�]��/@׌�OYZ��*L�8���[8���(H��[	0����&�Rɨ�/��p�T�ÞJ��s�����ج8�ѩ�N�!@�`k��F����,+����!��06�p}KH2�b�i��̷"�!��+�	�g�A������*]��^���n ��~fu��M���"�~��I=�Qvn����-��ضcq�-�]ԫ��|��=.�����Y9ҡܣA�wZ�
�C$Ȳ�=��W���!�֜�݂P��z:4r�僕��用���~�_�O��HiL����Ϋ����g���ì�X���G(b,�!<����ŵ5?	�-{�j��T�E�����9��vE b�8�޾��d�b����g97wU�k�9dK��stB2��ko��H�ޠ��i�RQ ��@�{�QKt�"�?`a�kX�����h�&h4La�EY�1���A�qE`���Xh�5�_;<�ю�/��gpΥ�^��)^@vX#�Wc��f(P�!'k��Ǘ�*�VŊ�a�����b):���Q�J�[}�3�4����� xsE�T�`�;��9�Uaj#��0&��$���j1�{�7�nb��,,�!ϰK�
����c(���U�8�[�6أ���2$xNi�ބ.Xv�q;i���W��)k� �؋I�~�f�0��_�/M�����&`��#*�T��ʟx�H�r���{�������В��S}��*��箅���y4�p���X����>K5Q̏dҬhAU�4n�U~��bz��I�	f�E6o&����j� ex��F�~8�̩�͓�����S�Μ��LuV��M�`�BmI��K�����nE��3���"ס@��JmZ�*����q?U�2Ǌ�#~�}wsW�>J�cޠ�y��Ya�B����}�×"L$rk��'ϲ�(�Q-��A��!�(��N���oB��GU�;�>ay&��S3Z@�o���'�,�c��X gh�Z9�~E�+�G8�z7
K��)B���k�DlU���"�"�9m�)�:�qp���8��� ]�(���/�,ߵjF���w�x�Gc�'M�f������A>�T ް���l�˂�2r�̊Kz���i'�N��\L���<�smI_���"8z�t�x�HnC�}J���bZ!BN��Z���ڕ%�`���W-޲nE�S�Yf��~P�i��*���v#��� �����4J������D���O�T��V\Ps"Գ�����ey>�?0���n��tm�ۤ�G�&JX��g�%�%sB�+X�{:��9�j�2���0�bF\���o��'��QH|��M���oS�1i!C���D��r[�aa">�uފ�����q�/c�$�(2H�RM������	���Yt�����
���"��Un4-Y~]�l��\��.�L��1}tN2��k�؆�����m�Ѷ�n���:uKdSkEJY��]�!]M�7"R	B�1J��N����Ŀ����d��S=�Kε�?�|��x+H��`L���1J���tKS��[AA@��΍8�9���k�|��:22�Ww �~��N t�4Xρ���'�}f-�����&Z��~'@�:��ۅc��R���!�;��)T�^�r7w�G���r_��-/<F�'d5+)����y�j�K���cB1�ꚹj�= ��VӇ�'�e�\uS{��	d��,���wn�S�nzID`H��RM��.�YáF(ñ�(�|]0�DY��KNz�&�I��E�l@B�V�Z�)�� ����G���6vuXah>��qGQ;��cDv�RYs3�����0���d�3���I����@�C�z1C�G�xV�n��責,�;���+�E�]�HdA���bD��p����νW/b��?�v�Z�.��a��qrF��1Oܽ�45�JTOF��o������f�q�Ę���K,-� LD>is��W��o�;_hB���2)�ۥJ\,���2,K�%Č�RO�yZ�bj-*�(º�!�"����f�;&�SBh�+'�[k^�q��/"7���U���Z4n�)��T[m����b�K��!Zv�$5��Ja��7o���_X"N������ ?��^'"��|�p;�ro�\���3 z�)��؉yN{��$�*��x]s��6�셚���L͒�w.��v5d��e�bM�'qpI�+8У�/���E��)S ��v���Ӆ���7�p�^q{� <P�9ɧ���ĄgsV�\��T�l`����}��Y������K���Z���%�&$l�
����XmVb+rpd|�x�A�Y��#��а��`���� ���"!"�ێ�1>�i�8ѷv�|�t���*��G���V���/]�~8�j������u\��#V �!��(p��LA�x�[R�ֳ4���(HyIA�� ��h�ۻ��A�~���� �z餶�&7��l�w�.e�ުw�~8E���*��#��6��H�(;0[�}bz_Z�s�������u�:��s��s��t��ت<�OQ��*+�?;S2��Hn��p$93��e͡����OF�?�O���|xy����<�CA�m^X/D�k�����1�"������\D�������h1w�ee��� ��Į��k�B�;�!�9�k���f�N��~Z���sf�!�*�l8Rb��՗V�u3�r�����!W��y!�54�UߕF�q"F���s,Y�bT�[>6��(E�*+s3�QG���j{���Ӭ%��g�������柚�K*�n��s�ѳ�yRʣB���C�g�"��[�jd�[��՟;]\�/���:�ьL���D&%79�B������TM�9a!+c��wd���O�k��^�+�O��	�V�V�2a�6!k#_�:�UJ2��3]��?ʌ̣iYSڗ 0B	ĴA2��m�����W;r{�"�Qn��B�����R[��b10 �pM?���L�ʴ�f�.T���e�sK��;e�����Y�G�f0�=Oi� �QYP͈���q�	#�"��P�	n��`�����g��k�G�7�ȩ������%2�i>��ړU�NQ>��������y�x��sM09n�N`�svúN��G�4�D����J�r����H�fo�D<hUM��3�)�-�B`9R���I��[Q�����]y�޿�GY���Fݲ8���C[.���"��O�S�H��_�S��H�ZKy�f�d�,�fo���}w�ǐ%}�෕v2�UG݄�`1�����:����~��*]���ڕ>���ֶ�r�?�����2k �d�J�� u9(۝��m�?�1u��� ��A4|�x��������(�>��τ�Tʆ�䑇�*�b��].���X���F6յy@G����/��$#!��s��}P:�e;,��L��tӧ2W���X�_ml(���r~�QLd|?�S܎�n��W�i���X��4!m�������8�׆;��כ����{�U]�cfK����lM8��	�?O���V���+��uz*�6�#,3��>ؐ|���:���p��D�����[K_��t��ᦔYF���R� I���;��2,�)���$YJ5�I�ۛ��˯lx>�s^�s�Z�#`-�q�G뎔I���<�ol��2G�]�d�
4������B�bK��d���wD]b6���7�4g�LZ��hp=����]�>�Q����W�@{�O���=��O_�� �cO�.��Ćt>	,V�s�5_�L]ެ��E�p��[�`Վ��]1���%����DoU60�^,ߕ�a����ojX-��:��5�Jm�t�w���SL��������Sxo%�����lt�dh���"��+h�"��≶Y(t6���, |n�н:��0��Y�u�r`�zr�%��#�7�*�ooZt�DOd�M������H;�&�0cOǠ�=�]C����ʔwӼ1�(]��K �� rs\��N����O#��z��]�`�qZ�����o�A��tf}UPc���ܬ��i_���,��z�Q=��rׂ��~����XJ�kG_؂}3A���4�� �
]R��-\�e�A��u�.î+��;{F��/�ZY>.VQ����ך��?jWW�A:��J�M�ή�{����m��v�b?�e��6x��S��h�aw�$Sgxࢵ	߶�a�Ő���7�ΛIt��XgI�5m0��l�|�,� \�i����N!�YL���&"�W=�o�"☁���7M6`���Pü8`^���U�B��d��)Xp,!AI_XT	PĒq�稑��l�J]m���۝�όE �������~�?V%Uʵ�@DP��~1�'�{����`����ge������� �y�,^W�Q��'i��T)4�� (���-u���E޶ԩ�;8��� �HUe�ڒ��*[,��Yހd���T���i\�-�%���G��L�6ϔa���|UG�cp�"]]�W���6�s����w�id+e�dL�����z�-�E������mnE�E����]*�y�~6Bb��`7����ݠ3"�,���	�}�{2��4-^L��d�Ҁx���4���J�m�1�[(�c�ٍ�,�vsy ��XU�WGRt��h��b��&���	E��\xr���e���8�T�&��H�v�"�Ы�o�˨���֏��Q����D)���9ӭ��]߅��/�{�g�nW7ֿ~m��9�S��
p���P���}IH�c�������sy_0i�<!��yː��ӛa�L�:o���~���;���8�]��9���;%W����h�3ρE�L��T�A/���d��-3�=�,�:�����~�Z�y��t�$X�1��cS�!�U���iZ�`2G���mr��jݨ�!�~��B�@د>��M"�������g�Y���h|��.�f�')�q��\�GڐfER��y�/�7��d���iŋX��$	K&AQ`���K�s�߈�2?���ү6�����`2�V��?�������`��}@�%�*{O�nk#UV�e�X�Ʃ�/�Z�uD����6���m81M-��q�9��6��8G��m�'0xӶS(�GG"�����U�Ww����p�c T�9v�v�IbM>��
��O�J��E�:��)G� ���Z�A��#�`��|Vn��a���Y�-�&�D�肖���D�tAlk��f�������������몇!"�<�{C{2 �FsI_����$��o��|_xwbV�`E
� ���) �r��f3�-�X�WjK�T7C.�FRֆ"���7�.��e�x������ȝ��7�ļ�рE#��?��k����#J�?o� ��럤�7Q�ֳ�|��%�rޏ"x���;�*����z�ݑz�5���t��Avb�����*��m�`�ɎM� ��&�,B�Z�[%�7G���_IZ��J�k�.��=YT�> Q8������δ������w#�
b.pK=�G��;�/,հ�]w��C��d���?I���r9�Yۼ�W傕�-�G�33-	0N���e�Ni9=���%����'������o�I�����G稐W���,7-����ųa+Xo�|�3r�-����pn���]�Y�DT��k�t�ۅ�ʗߗ\xq�ɒ�8�A����Hc�A�pȾ�� ���0$����2���5`��N:c��Cv�����ҿ�O����k^�FN�
��f pQu�G�3 �q�P�z`��n��ry�A����ϳ-Ԧ��'�Tx#�	>FY�e7�?��k0W�!��K�V�@]���Eݲl��t3?ʛ֍��k�,aڠ�Y��r����n2�S�O��L�A���NR!A,K`i(�
3yxv�c؜����p"6yڦggqm4o���wTzJ<�у^��%�
Ş���v�n��e�i���k��� 8�wd6��h^91F�_��s�Q�|�d�$;�M%��`�aSſp�����2VB��ql���S�d�J�gg!���Y��C~{���l@�0T������w$��;��n�p@���"���߰���;e�r���A)̄�р١+��N/��-cK�Ժ׮w� ����{D�2ɶ�hp��.M�.��06�\�~��<���j��]C��D���C�^��ȱ�])��ov�ʸNpfe\���o��R\I�&��s������~���	��_�KzKA�IC����1�<�&� ��!��9�8�ې7c�ro�H���h�7Q������Ne�|�^�r�{��\��ⲋD��I1w^EA~Ag�ͼ�^60�F�ݜ$���呒�ʁQ�7ʽ����"�X-���k�;�H9�P*� ڝ�5I{�N��<�o��I !����������Q)��v�K_+r��i@�� ��jC�6�=և�#���>��:�4�D��p�s?�F�D���׷�P��w�c��Q�b=���9�ޅ_�_?.X�lÐ^��4�f��D�.e�%�)�/ܞRWH���wU��,�K�����b�[yE��~xx�o>?��j�\�R+� ����p��w�Aa*�I"�;leI��H·�nSMG��$F���,�P���!ā�h��M���lQPR6HI�E�15n�n�9�� 1���ɆGs��'�k��iH\u$����4y 7���ཏ_��*DM����kQ�z޷CjvX/���k�b�6Dp��۟�ʹF	��*V��B~�gm�:��9	��D;�<\,� �<;��涕}��IX,��&�5�RaG��́Vgs��cJz��D����i��'9����8�O?���|v���ٟ/�Ґ<�I���#u��F��G��4��ˣ��雚��V3�6B�3,u��.Z��s������r��B��8�H���<���q��S�o�t�¦�Q�9(���i��h�P
��*{Ey�`/R�u�:W���N��7S�O2ۄ�ޒ���<�dm������D��(�|���7#�1�v7�a�ȿ&��m�Jt2N�!�֝���(�R���Pq6r�fM�{y�xlu�u��6�p6Wwfj�B�K�"�yi���m~H
| ��k��h��Ww�	�5eyx�j�`�]�AN�b9��d�b
n)�,5eܞ�)�y���74����J��i~w1�?����\Pg�<�����Irq���R;e��9��@B����k�T�q��;�;}H.@��k���K�HЦ'��p���+-��M�(��8$�Ϸ�\�E�l��gH[~R�:�H���`�]�M��Z��n\gmlG������骞��v��[����#��C' B���Z[�]%�	���x���N�g^���R�u(Q�oe��^��=�3����9ߍ��;�J�$��xDQ�K���]��z+����T2��|�!6(��)�I������$h3dRz���*@Z��i�,$@ ��P��?C�l�L��xs*i�A�10��&N����_�^,~�ϖ�1Piz��T檦VG{�[+t�B0a���lHrP�X�i`F��|�R�p����vѱ�H���Z�N7b��LdJg�Qk2�e�^�ko������`>O�HН�G�K)��2�Ii��F:!��s�͕�<��#�6+٬��/v���@�f�鿝t���zz�����ޕ��2���F?-��!�n�2�)r�;
�g���������1�V:?X�?��n(�g;��OA��tT>�Fn�A�d6B� ���Vw�VH�1�>u��-�_I��y#�[�*��V����m�eB*�H�����Ƨ
C�al.9�	@
��wEgٹ�I���1B��/b�������b�*�^�_��"�9��x�~
���G�f���s�]{��K+a��D����X�-�@0ћ�4������=��".�meZ���ŭ�v��o��i���TU~z�;�"��b�su9w�GC��Ҝ��bwy�����%H��B��G��3��g��rG��S{�CQ�	�4�O����]�?^"����Tp�{����l����S}��¬d���� �Z�M�'���(�d� �]B���U������(F�9������n�7�|z�W�Kq'�.�i��}s����ӫ��	�af3��9/#ZOpU�T|�ν����*c��;��ŮNy{$w��5J�'v}�PT".��ܶ'��ES;�$�R���$s5���G�M���}ՃPf����@ ���i^�o�~W���DkMމd��������'O^i`7�]��HO���<�:�h�"J,��K���s��}Z��vd 3���<���z���R���7���N�1�~�m}�n6��v�W�5�_�вh=������Έ�L N��k�nw��q��e���N���2�So�y����:jJB�0������.at��<�����mEc�*	�\)i��hDʉ�����Y�[>k��*��?'���{��i�$��R�:;:n�v��� ����rdwR�����]9.�3�K�dƛ^4�[�;�)�{f�5mE5�#�����R�cz
��`�s-/L��AR6�:� ��Nƶ��@���j����I�C֌q��P��K0Ыv��!��+߾�T��}&��^ �Q`m174�Y�(4�ʯŞ1X�?ъn�KOL�/��%�	k���_����Y��=���f�TGO��Q�S,Ӌ��l�Ҡ}���֊6!xx���L1�!����_��#*��^�N )�E8�dt�!�����t8�Ibm���1�;�x-2�W>b����.Bk��x?eb4��X݌�zȗ�M2��Ta����כ���WN��o�ޱ���WcW]��"C_��m�!�]��ף����rؾ�Q�#7=��;��S���k>��?9��(�N#|b�qK�L?���SO��S��=@�p�_���~��h8(������K��KM{B���@��Y*�=�p/U��`]���� j��Ģx�V�����$!Ù��$^�ה���pPyY��f� �4aq���3�Icucm�'��`���I Ѽ�U��,n�z��B�;�	~�(�Mg��Kw�E�2!G�3` t+O�����K�с���<A:߄�F=�����`� =O1L���HO��	�|�ٜ+�5�/���k��l1MO-6�<�%����ݖ�(�'}͸�>�_�=�^eP�U2b�8�ϣ2{x��:�< XQ��i���i:�����*�3K�?�Eky��/33��5�)^���D�%5�(r�yo(;������xh�&�w���&meP9o�R	 � ���{.�uN��5/d,��@�Ø�E�zTrREjG��֏�>p*1��e�ܬ:�c�����R�\��`#LJn	-�P6y����@a��7�����E�	�%'�k��:����e�p�F�Bm=������Yѕgd�*�8i��p�q�0ݶ5���vP'k�h�>E�X�)-��\Rlj_��NCs���1f@�Tϖ�8׭��u��F���1 Rj�x�����+�Ğ4���'<�!q��er�Ǟy����!L�//w �l�^bk���˘�i�T���Sb����t����6�e��<E���m�G��%|���}zqu�/�n.ޜ@�Q8����H#Ҝ��i�o?-k�0�;v'M�d:�z?��B�k.�o�9��4��t�x%	B�(��'T&�)�W���.�<����zH�ٴ�ѹ�PV�p�K+��� �<6n5
2)w�t+���g��k*U�{*�?Cbūs`o�!x�V{~c��Z���!�M��XU�c�����vG��I��3��a�d����ڈ��YH�2�mF����f&�$E�{�h�����60"���ζ�qnK�w����-�63�lÅ��%���:@I�)5�P;zo����L�.��Pr�U=3��yiL2���b�.cI��Y���1s��X+�g�U*E%�N'�\��(�;�ËH�|�ћ�ea� ���2�����_\@&���+�{�]b z^� �Z��f5�S&�<�=�y�Q�|O�IW����R?Od4�m�ƞ�erM��CR��ELv{(��-vp2�=f�1�#T���`�ww����ۜB����L�Q����E�"�*\2�g4t�9[�O��(�&�[����c��������a�
�
��n`?S��qL���=�2��b�󫊄z�C��*�*i��L�MWV�����ڎ����̊|d����*��,?�1�N����o���6�0O�z��m:�`u �XN�n,i���b�U���r����<��U�$����ZD�����V�n�j��K~0W.��p��:3ȸ�#�,��3ߟ���/�b���(Z�a/F�\�b;b���9�������,��-b��D�W@��*��~�I�)�T��5,k�R�5(\)Y�љFE0׵2���о9��BQ��-�����rx~UvR��΢�la���E(��*jl�G�ͣ����{�CzmAB0$�4��t�lf?}������0�R|'�m'D ���s��K�Y��3�<?5>��֋������A:�}FP�!��?c^�_R���H��v���o}��s�����������\μ�g�oI5hV�C�������ۖ����S>?zC�M���noԴ����b_�vAƼ��6F����`ߙ�����
�C'���َa[+7g?j��*=>6�2��~&v��@��U|�劉��T�@�S�܄�	)>���@f����"��q�pgd��>��G̚ޓ�.(���[1�-��}v���({�B��U�ǝ�B��J����'[������5?��{�;o\�K̢k��8#���v�_��i��;Q�)gy�P��Yݘ��ē��tY���.?���3O���Z6a�f8�_�ڮ��##�&�T���^3}��+K���iϘa����w0�|�ܻ? ���=a��BNk�u.�*D`
l�p�@	���]1�7TC��7jߞ��y�}�1�uv9�V�/ lȚ9�r�߀Ů����ߘ��=
)��!���3y���ˀ2W87��F��s��H�j�)DrH�/2c@��TTE<q���q�n}[BW���;��\�.�b/��+��S�?���Y��0���R;X�(��a	���Dy�����H����:A-������]�&����Rw+��K�p�p�*�h���vt���%^�eWV���Ż܌�Q��o��s_�X��s��ܛ6��˕[T�89��|�a��W�����fP�y"j�E�TmpĜ��N���K���� �I���}ar>��gi(o��O�5ܴ�f���i�q�f6��	�X���;�_)	���@��BM�Z����;��}��?C�0���[�H�٧-�'��vi�{���`���0J^�����#����h8o�%ޚ��7��ݳg��T(�Ήzg^0�D�
��Yވ������l���1�㼶;�[�1����QMX�"hD޺�ׅ[��N�s��^�8�O��F�B�v��S�H��vJ�Ĺ��-*�L��f�-F�1�l��s��
8�x�}a��!����q���u|A?�L�VͿw�u��},(��\����+�A'+�-�ū+���U_�b�2��c�w�7	7�Tv~�Bq��VA��W������b�E|I�����0-3�͛D!���ńa���F��My,/������p]��ٲ_�E�J��Yȯ�������!����^�V��l�Dt��G��A��Ys}�l+�|:%N��_�����7��I�dW�y�j��5�a�,ᱟ���#v	�i	ˤ��[�ب���A�M�,��(M�r�H�J�$���j�z5
�r5��g		���p]D�E����<C=O�F���k:6 �#�5Z���I�u3S�o3O��F�.�9UnF{<'ހ�a��2���a5�z�M&�L�^�`�ۥ���+ż�f˗�\3�-���S�[�2Q��Z�Ci��6���Q)(�h`����F�c�����Vv`!�j�K�����o3H/��+it����ڞA�1�j֘�*�k���+��n��;�T��	�$�(ʯ7�*kS�]�-�������5(j�jL,���G��`A�T8O�J9�͌������>W��� CZ]N���p)�/L�H�u��ymE���"�aIlh�,'rܛ��9��&��khL�\�}s��.4oe�]�F�'?���/�Y�z�z�bC�M�/�+���iu��^A��n˲*�B���o-���sa2��]�Ă��8tr��G�	[\ݞ ��.��F~4�3v�E�\��dW�/ �
e�PU��L@i����G�T���@�éDL�[[��0"�؍�i�C���)k,�y�|mC�à�(R���P�l+�9�?��7�`�Q����{L�/�WU�Z� ���Mm�#pr��V{�QW�������G����wB����"�l�,�	��dc�տ����!��m��|���-̹R������ω��B>Q�cmt��1����;U&ٝP���z8J���ʞt*���sU�ā����k�ɔ�9�]�}_��Ǒ{$�+��U)�1pT$!c��3���c)�mv���7C�6K��v����d���FmcH����]��?�M�m,].E(�ZQ��
ͼݻ�ӳ/�����j����w�
$��{�� ���|��_s_F�m��7��
*.���'��@�Q�Êu��<��}��r����
�/c�{�+Hz�i	UnDdH s%���eBf7�D��Ӷn�zX8Wgm{�s����x�Q�.���K�=a\���J�ܿʷim[��R�M�e�<���B��al�
{�P�O�tV�j���� ��	����|�qfK�bo�P� ��s�(p���M���QUdu� ��Ż���I^��Yo���q�$��Xe�b�P�H�[T�-ԡ,�.����g2}��P�2�) �*i��^Q�na/��~��o(H�Y4���u�3R��FϨ��CD	���#2��2��{&;���Zv�-��RhZ���3"(g�LӬ� ���:4�nZ��Hut�c/ܖ-�TB��k���q�ЛR1���-r��~�u�-��;�de�10��>��lc����e
��z�,J��\�=����;�~D�����b^E3�d���2'ÎL5|���'8���:����ϼ�\�v|�#�3.����
��WOJ�ٕd�F#�8ښH��e�G�)��,��g�Pɺ~��i���O����x�L�D�(�v���1�&�5�.�n��x"^�= [����*��� 8;?�2��ٝ��[m�$���� �j0^1��be��À]��b%���*���2f\��pLV�(a-"��yêd7����C11�7E�g�+}��G!���o?�A�s�bX��a-�fuB���Ă�6�C��8n�Ϻ��BtS�^��Xl.}��r����7.�h���Q�/�PhZ�4�#�u��C�}��i�ӓw��5�?^��6�~��J�a�q���@( go��҇$�<u�7=aU`�i�[ٴ�߂fx�iK <_޽��8����U1���"Ν�r���l�`�۲�tCӂ�j�B�u��8N�;������1��h�hC���"�����!�/�^(�~5���A�j��f�f=G��U_�g�r�VԦ���f�F�x�ZB/���<�D�J��AbQ�>)�uM���A� Nr�3ph�P`;�
��!�`\������QU�S>���Gl����f���W�?,l�//x�J09;�Ez��;+�E�����i��/���J�����@�Y��&�IU#�y|�M�ٹ�S,���k��bX\hD�NL��A��%�^�a�6�ɽ��̀a|��ݯz6�P���X�d��`�� ��3]�{o���/u�2��u�oCfM��hL�}����w�Id(�rZ����wacŭ@�oP�����v�Q/����BkыGDlwvj��AP��s�*���h$V�������	������$/��ı>���x>�|l|�~;���_z��4�%���w{\�V�� d�X�D�}�r��ƈ>���3q\H�ˍO��Cb6i�sp��3fd
��V�J���ow��&<j�C�S/d��).�*@TÒ)���-�=���,���nٹ����π��No�|8V���.��j�c=�S�;:�Ahb�Y���h���İ,�xf��X�q��^�D��n\�z����(�r�0Z�!\tq;�����FA�)���5�������b�{�-�C繿F�n�:Z���A־� �X���G��pҒ��<��J�m�ʜH�������q6=Zɑu�A�S���Wvl� �f��eZ��`����I�����ap�FP#A
Q���_�և18�s�\=Y�l6��X�mxT�a�A@偃P/������vg�؟7���u�t�� #O�e�dnQ�tgb�R#r�d�,:N��cW*��n��,L��F�#U�2���W/��Wdy���M����d �כh��Nk�r=�p�1G�7�3֮ö]T�G(��jM�d�y��џ}�'�+�1�� ,w��/f���BXa��3��,z4� U$�������Yg����D<��SG�Qpt�'Z�ᩕݳ5�۫�#������R�?���P����ĈS�|�X�vUn�{��Ȕå���0(=�)8�0�..*�G����?Y�j{�􍭀C��2f��MR����5lJ)�2�
�`kTs�1X~�z!P揵���z�<��wC&sP
>�ך�{���O�ṏ�ج���^}A%A)YL�wE��'K��W���	5[��m��N3W^o�m�T�f	*�\a���1}S,�K7���Yd��S~`�1����VbGS�fߝ��*2C��m:��o����YzW��ݓ�*lL�'��TБ�2A `�s{+7�F��%0�v=�5
��������"Z��Թ*���A������i�^ڎ@z{����:.0�d�g�B�#3�xv9N�o��i�eMR=D�
�H6Jo��sS��.h��ǣ�̭��%���0lIP�5J����E����=)o?o�핆Gw��d ���?KN�(�6�GˣY~�׈�����vO�Y�H���c*W-L���LY�~zh�?p���@c��hE������D1)w�ݛ������zۯ1�5���&n�ȇ*�z���4C*`���&�ـ"!pl"s]^�
 3È�rm��I��
ԕ��� R���-|�?�su[<ayU�l��?�@�����m'1�>�c����U p����y>��d�l�q���2�K��#��3�n�U�+W� ���&�j��ǡp�q��w���������=��'��̨�����Y��Q[��� �������4����G`���v��5��g�锩�K�ΐvN�[��9�n�a��&0�7	T%5o�ҋ����G�2E�?6�ư#���0 @���mT0�<��a�������臏�G�POL�3v�J���]ND�T�p�	��|[g�0t��0�
/m��s�.T�����o��ՠG*��V`{�/��Tͳ$��\nt�#Δ)au��+̧Tvo�]	�,ŋv4��K�gfx0��US�e��������B,(R����FgO�x�9���E�<>���qud��;R�Z�QY�K�����{�5��#�|2`7�<.<���VB=���כ�ݍ�[�!a���|�^G�w�����`.�ŉ��@mx�T?�s�r_�����N�v� ��/Y˲�uu�6I�7�#��G#LEӴ���6���*O�gK�Y45�"(:l}]��rLƱ?�<n_��Gr�ɯ��
��} eI��VU�v[�</lg��tT�
���p�$,�,P���:�����[��΋��0n���m�m�i�X2�V:ERg,d���~�/�ڟ�"�DG�&'���5���a� 5wӝ@�AJ�Aly���
_�;�-ڬ����6CbzX�/�2+r�GZ��q�.E�X
SM��Ω�2ɪ�ZiR�H��	!���뷴�,<Ӳx�����3�
k�ֱ�EZ�k6Ś
)��L.mt�tvٯ���H��{Gl�0�E�i6L#^�z���IKT�6��>��w��=+��5Iĺ������O(i�!����W��_^V�tؓI`�=�w�f9|�O:)I��,�T����鋯'��$�s�ϚL�
Kzq>q�묂Q�Q���Dsπ����+�"���8��A)���u&�&L�õC��� ��:�˶��ܫ����}6]*K�A��"4�_��x����0��J�	(ҲKdX�p�����S|�N�?�c�p���1�qnEy��^��a�n�g�P>��/�&�/����ǒ���Z2n�_hH��3o�%�u2�:�/�g}�{H�l�0"�W*��v�l�a�����28�0��e�uZM����8I>�J��t�.��^�
V3Y�[�%��a�|�m�%��k/�`�0q�5\��d��k���2�d:b4���a.�1�!f�#;U��_�]H�B�R�+�+Lx��_e��Y5�i5}u:`��n%nHh�y���@�����ʱ�f�Ś�`J���{G
L7�=Q��s��e����ߺ� (�����H3b�F��$���Tm�fk������c<~ɡ�����	5IvY����t�T�dam����-�����|�����Sњ���8�m7�t�F/�	VNy�H2�ef�˂$�#�2�6���69���6[���.=ԍ��Ѩ��rHN9��H/�������,UK܅e���"�Eg�5���t����(��eɮ��:�݅7G�MϞV��l[u�xI��1P����QȘ���x%gC�3	X?Z���ҵ3�F0 ���Ō�����󴲳U��p��m�D^yXg���Ac3�7��[=���!�C��8���IB��?��/G�W:FGX����S��ע�*1�£t����9Ár�~[�s �[���t�vG�+個s�q8|�GE[{j� ;Z�>TM�A��\Q���m}WTt��|D�d�8��*� op��q.6N���/Q�S>�j����"/m�z��?����@�����$���p��h�t�\����r
b�q<\�.]3��S�r�J�� �$�P$l�z�&hWdQ�S0�^,��i	8�u��#�2�7%j�� ��0>k?N�wT�n�,�x�T��a8�S�Wvb��)ٝΒ�tw��S9��>��ۇ�>����:$���+��[�w�L�=���&-�O�Y�pz)������Ťc����.P| �A�
���� M'uSB���JK��r��mI�u�4۰�YP K���
܂�_Ԡ\Ox9OTg�I=99�J��ݍk}�A�D�)W�K�_Y*�b&�r�����ȵf����%z����=w��(�m�"
���h�N+.FS�`a�����d�X9U��kg��@��{d����H��e$�|��]�P�"rR,�:�8:���)- ������O~_IX�r������ּ_��fU����3�G�(�I��YDW-�
%�pJ����Y�0����R�y�0�"^~i��Ӣ��W���mN��sq8`�Y`�X�Q�C����z=�G�������3p��_��Z��u��5��ڜj}����$y�	�&���P>!�$&�Bƀ1�^�	2Jz���ed%%l�}�+
w�A���g$A��bz���yt<�)������u��=W{�t19ER)�]S��8��ľ��j2O�hk�=I�>�c[�!X�8ցEl�k�s[�`0;��<��	��H!C�X�oݞ�!�.h�`,�~7N��:KR�P/�Ϸ�^�>b�zIIuY�O32��JYf��Q1���P4�t�>]��kQn�]�yW�-�����p�������61Rk�kd�K,�����VPS'���Q�pS$g�՜��:s*�~���seN��n��f�ܟ53|+���V��2D�C'/��i��3ơ��(�i�E��Mu[Ы�L��UFDX�F&�Ձ�KJ	N���!=S�CcZm�?�>�S�d�t��M�W�I���-~���v�G^�j'�aI+��'{W:��Gx�6�6[T�})�(�r:=����U����T)�l_#��:�����tf��r�G�d�)�M����
�Ku�la����ܛ��6A'LФw�;lʮ�(Z]n���r�A<��Y��$}��H�T�󒥉�q�Ÿ�_X3���34�=��p7�9�3|��lS9��BöuՀM�z��	�v>`Qx5^ȝM@���7Os�6.�E��-v9{,�J���Wυ���Ę���{�i9��G���@����v������+��2�)�k-F������������By?�-�I�!��FGH���r��U5���*�a�o��<�����w�{|Ý�� Vlݺ��5
���5�h=m~7g��*W���Q)4����H��jTt'��J�3^Q���]� ���S݀Jq��j�U?��c���!
O\�zm^�# �:)�L�D��7C��DC�z(�;;�_L"�����e࿍3��e�e�s�@�~�`w�w�1����$��h���=��x�۹��5n�kWft1;��2��y? �|��:n�����V�t+��|#or�L�+��(�𘐎R��%��$M��yV�.�c��T\�zE?��'��0��%I��倿���
��K!�q��6X����P@ٛ����w~��j6�T�+����}�V�T�\��H-�t��2�+�\�h��-�
�&�#T�AZhքW�Roۘ���S��[���|�@l17������`�	L���4M�@	�z�Yp��5�<.�W�F����}��XV�����<,�o{C*K8 N�/H�L�C ]�غ�'-��I��ِ�@�,�$����csm��;R�����'[�� �[o�$��j�W��Ռ�̋d��V_����4ļ.�[�@�$�/�ݵ��T�/5S�˄��?���t�*a����ӈ�9��DP�<�?]J�Q�Ùٽ��(��х��񍠳+�Oe�|�x� ������ScvS�pRֱ{7Z^ag���>=��$Pb��ȟ���Z��U߃�Y����'"�������6V�(�W��s]ϛ�%N�mO\�"��]� y6Fv(@Yr
kEβ}���Ա\��G-�>G�-� �f�o���E։!�/�l�UX���e����in��d��(ԧ**��1*'	{8�g��@��a���z�_�v��k����
|��3bP�G���*�y�����[)tẠ�k��A%C�V�)���a_#9��F3�h5�E&�.=�ߘA�k���u5�J�|�K7nd�x�E�x4ap���}0 �)`�V3�n?�]�]��b�Օ8Q� ��ʄdxƧ�N�q�!���O"A���(�t���o�?���Au���-{�NӅ�\��lNS!��f�׳�>��O��Μ.�����Ǌ�sM
P�윌��Kؼ�����$%���C���@���v3�$�f�m=S�
�w3/��bm<j/_Nk�������װ�Ytxl;O9��Jە-G��F*�T��3R��RH6|hwc�$��,`��yI()��9ġ4�9�4��mVM���鳳�'�G;�rQLmO=�+k�y�x���g�j�>�{�[��]�/xE�E��hf��ʮw��4��EU�Z�xʞc#��[J"z"j|\�oֲ/F���=��"�#B�����1}4�k�N~S�Zp��T�1����ܦt���$(>&"X�+���߷�������V�HPKf� g��YiL�	�$oX�*�`iSôL�q,y�	uPm�W!*5x�������E�靳����X��vو:R	C�G�ѐ>��@�~ '୙K�Bx~������+�V2),�?h�"N�f紺������K�}G�)�h�7�� �t��E�/��*{L�US7B��~Sj��\r�fVd������8���]r�9GEln�M��������+�F��g�j��Y����몶ŧaF�zϛ���B�;0U����mѴ���f��h��W%���� v���vh�+���>�A x�tG��9j�7�d�I,sG�
��nW�p��ߒ�DƤ�A+)!�;e��k-k/��	3d�v�?`�d�<Àn���r�����i�+�%�?�E�D�i��Xh�� ��vH·#䩥�ހEQq* �q n�R�U�!�y[=��/�G�/���ζ� &����4�,�`��ߴ'*�7ST+`��[5 S}��M)y�]'T��@%[�9Sk,�ā?S���>��7�h��#��D�%�tcHZG�qk9I")m�Kvg�Q���@�#��S����ʣO%݀|f���oV�E��ҷ�.��F�LW���x]?,ۇ.��=��'!��|�B�3�!����h[g����$�Dv�Y��VG%Rԗ����%^���؏�%���[Ȗ1A^��9:���Fa�'"*�'A6V���#u[���0W�-��4�K�b0�
'�N�I�~ZK���5u(uP�L�D��lOf�l��V��F6�ָ�ZR�� �x��uk�����Ǉc�I=��6.��s��UQ\΢���vB�4�4�(M��o���UPH$�������Fd�g�w)W�!�=܋(X�-O����P�Z-θ�?r�㔢)�X2�0Ç�Zp�����+���#�$�΅	�E�:f�	�'���/��_m�~6Ӄ*W:���s�i�����԰���X���7�K@����&� �V��d8�wI)���'S��7W���q�8i��m�`���>l�釉������A��F�j�l9,R�-&�+����r���d1�+{�֯f�o�5�/���$���Pb�o$��'p6�^��M�%ovP*����N����]�rL����-��^1I,��)�	z��v`�Ls4ŭn�DJg���ՙk�>D��2z�
~��%<q���W��֔��!e������}���T&>>�i�$.;0�R⪠[1�x��P���1a�r`�c��,}q�h͋d����:Ÿ�qF�<��
>4�G.－Y��F��w�S��!��(��,#|�~Ҙ�/��ڕ	^����w���B?�'���pO]UW�4��]�)i�G��I�F�zi2ֶ#qR�Nk~h�^KY�+T"-*՞5�n�^�6�vH��]w���������Dl"{g��fi�[�K�� #Xx�cY��U�"�Z�O�+ޝ�G�**@�O�����%�i�y��A �e7K�������:w���z\6GԱ�q|X)�N��=vu�>\��,8@ɲ��ϜPX@��"Ӓʄ������ء�в��B��2=KܼƠbH���#?��酜�	w���Dy��]پb��|2,�i�.�͖Ȍ�����:~��%3~ϟ��4�����r���%�am�DK�#�z���\/bJ�57IF���J�N�4��Mƙa�I#�����V�#�
�¯�e��ֽ⊭p���<�h>ا��kG��
/��7I1��R,�*(���b��j*�gZ�p�a�gS��A��k7>H�yvֶ>?ɥ��ĕk�CsT\����7���$�R ?���갹F��Fq�nįg���>R?����S!�����v�k������ݩ�o[�_v�yw����X\u�J!J@}�?��S�uM|�oz���wY @�|vV��W��Ӽ�=���%��$(��Ԝ�T�I�[h6�''7�b$�:�3��Ob��t�6%1�{E��J��^&�ˮ�d ,��� �^�w�.��
���;R�<�����B�'�-#�˿iS5a�j��9��I�w7 �� l���X(3*��j�B��*b�x<d�Ed��� �5V#n�3 WUԫJ.���rX��p>��I��J��_#�MO^l�t��D$�Z�M���9�"��!�/�D�����p�Ny�: �
��DܟŃ����j�����jȪ��yyG�T��$m/�(�҂�T{�;N��}�C^A�ɄB�L�{����~����ٞ�w��ؿVC����uk�wA��p��}���q|:JQVyw�1䮢(P7�Ś����B���-]p�,�����˳QZI�a�p]��u�Y�̩(�`����>�*��*vT��(���y\���P\���=�F�m�/� �=���u=>_{��V�ݙ���h��G�Xs!��_��F��8E�M��9���c�f
+<Ω�WF�.\�i��.�FLr��5��@�
��ѓ�5?4���K�3� ��QXM*�����H 缉`�����3�0�5��`{�>�p���2S��������T(����1K�H!t�Ԛ]��&��a.�K(�K�8�хNH�^d�8�3�4�g�tDOX�$/V�A���$ez:ֶ�s��Ǚ�>��>b�
ι1��ѐ����a�'�z��)��S���0�^c[�~�p���M�Jt�ܫ�WY���L&al����d���nJLg��s��ð>6���ލ�z��b��� 	�Q��G���~����E544%H��wȣ�m�%3�$EO�A�ܮm�)>C��\�A���z��J��L��Mx��x���7�rhͳ䄬'� ���a�#O�Te�u �>@�S�[Nʜ�}E��X�Z	��N�������~��+��NrG`Pfy����:���뛼�G��� ����i�X���ҍ���O���8H�PD;:�(iMTѭǂ������ſ���p�jv^�i+�{Y?�ʽ�&��xE=����ę_� ��A��p;/�E��v/�1���6j�ӈ�mY�~m�O�Ux��1,޺���^uf�Okㅳ��F��U]�mA��:9#E_h�)��� %7e��p{��<�Q�Wɼ��C��A���������(_����m7�r ��� \�0r�H0aE��;���!v�+wO����Z���}k�$F�<�+���� F�Qf�0b���	�ڀ� �m2�=�IZ�����k�)�1���?)�e�#Z��a�s)���GXu}��v,����ͬ[ya�.)�'m��&���K� m'8�P���j4zp����n��ؕ��>�m��yn��	��D��-�9�,I��y������D�<���ۄ[�>8!]IJv��
K���+���o�jt)~�B���1���jD�ڐe�Co����Y]#����Vo�Va7:K�ٟx�Z&�~Xj�K���yxV��8M���ysKIpVc��
*7BIѵ8��_b����a�A��;K�@Z�C�pE ���ke`�'B�\v��y�9��e�7���s���S��ԅ<GU[������.�$ȗ���=��g�C�Z�C<��8=�+Ul˸��B��v"����M�Ҭ����'�g�Ĵە"rZ�V��˖�um�-�*�:�v�� �v.P���E�7����q�%w)9�<:�6$��t[�,yR�V��BJ-,���������b l�8rN�`�W4�.,PA�&��o�AXD@��އ}�1���f�� �A���Fw�	���T�����B)h�q��Ʈ�ÉA�
,E A�Vv��b����,m�Y�[l�.�PN�����"�� �����d�W���S��qԌ��c�W��p(��Nʎ��u�&�Ƹ��RHBdɹ��*��!��Oo-/���]�ֳ��4�g���Q�����MuD>�@In��{9�<hDQr�Y)�ס>�x4f.:B(<�0�O	����X@�G=�q�G��^�ܙR;��0"3���>��o�����6�����1���ުA���K\كq�]Ca�f9k�nQ	yD�Ş��%����)*
�slۈ���3=s��Mq� �|����r�-ۡS�IO"ٌuL6����p����/f�@�!9 Z�kE{{�#U�XddA36l�e���r�)���I�<�qY~%�O}�R��a*�mu��ڄ��<ۭ�ο<�����l�
�p5�r�L>��k��~(kQ/p�(����d��#Y+� l=�rW{�!߼�%[$3��'�}���1���.�g��u�|d��P������DcH QU���Z{�bP }��3�v6���E�yK�쥀�qP��l������	�%(�n���4y��"��{���U�ٞ%�8���!��'�j�x}Ũ�F�6GD���SB��ʰ�»�%V�R�X
�w-��.��Nsa=v%{�Δ�WR�.R�|:K@���s ��Ws�_�ӧ�� Ε�D�8��h-8�S�q�I ��)��$��S�xjX0�֎&<�zW�=��W,��F��=�X$a�/FNj������Q���_����SP%��K�n/��|`P,�ٌ��e�=.���������c����MQ��_�kPy^���U�)�mEb�����V+=*�i�7u��h�H���.zC\3��,����+u�`�������&��܍�`#��:|3���t�.�0!#���v��B���.����A�g�ъ�1�+{�0��$]}ϖ��f��~H9ܱ���BS�!�h�e|�����[�~��Bi��,�q�c�hV"�~�p4�A�����V�pi��	A �Ӣ���Ǥ'���E��L4�rc��B4RD���GT.��+�m����R�ec|�+��8~2�QSy���
�Ϋ�м�hRB��En8��3:IP��\�<���$�Yƛ����
�C�@O���-9V޸'��7	� Oϫ:NPZ��&(3O�ز��/|�~�=I'�Ե����.��г��ů7/�7X,W���)�"17��M��Zǥ7��%�U�D�w_�]��#7$�hnb�(�<��r�tS�0��i�t�2�}��_Ɗ�p���&�L��:�uGm5��Bi����/6���h��:쳿�����[�@���g<�u��J�� �t!Vz��zM��c>0�80�,k�1!�y�O�ҭ���\��H�`��W�Jw��M�Q~BJ2����\���y���L���@BQ���`�/����WOz�J�!5�F}6�
4�v�fK.�cn˩%";cl���9���o�^;�X����Mǳ��H0/�eT:L�m|35��-�W1�OA� �D{��Ɔ��ٸ<�k�=.9F�D*�f��z�#�Րܪ�R�;J\W���uY~a �(0��7K��V>)��gs�ɜ8�."\���UΖ���`iX`#�����Qʖk��P�5#����zj�%��у�F�_l����=�M^$̱��DR~|{֋X�%�T{sQf��t�*�����ĽЩ�v-]B4b�!�F	���%S�9[i��EYe��i��1%@	�jl��lf�Nd�B��4�����ASQA���~~�ʴ�v�p�#���}Xݤ����9�9��n禞s��eE�!ͅ��D�;p,�2c˾�����G�U���VhZ��¼�m�h_�j��3��	%���r?j"��w���m�'����h�����QWV�\E�������LQ2M*.�uO����?�ֆ/�����0S�yh�#*J.Pm⊴bj`�����2S )���<_B�����/Q�e��3�gA(��"�qd�� G�\!��i��w�[��	�4�u���K3���5������@џ�@�NK��%Z�!�S��;��w�vtv�=��"�_	���B��������b�.��>_�� �'qa ֯��@+i�;1��q��б1��D��#�<}m�����P��T4AO7	�6!�ϵ�-�K5++[ЫgW��h)��
 �I���)9>�/{U��`w�4�ɳ����4�^0[U9�s=��p�]��tL|�A<��2����4S��.'�/�*B�'| .z�|�:"Ü%	�6o�@�5{X�W��������V�� �u�EG�7"���3�HFk&nt��5�\�2a��q::��w�Fx�ߜ[z�l���xH�喥���y�gH��	�9�%��M��y��߀sS�{�8��2St'n���B/]�L�޺���@��3;Cu)wY�^�vͤ,�k}���SP����X���@�<6yq��ڒc��p�Okw"}E�3� �� �p�Y�>�_&��h�79��R5|{67HJ� ����+��D(��vU��� ���FFsil̻u�%�׵&�2~"�6}N�9&��\��!�(P����04�06k��S:%��~8+l�kP��<$V�wJ��S��� �JX��f�(\?���%��3� C�3���������q� ~۔kND��m����n*?�Ѹ�I�~G�&��	�z�r</_Y��+x(�\- OŒ&�'fX�9oa��Rz[a_���(R��I��@���a�a 1F�&I�9��zg8=���c&�)f��l�.���E�pN���d�������=�"��O��.!��&��i�K'u�MR���us����uEs?�|��2�Ñ����S0��� g�w��6�m�X^�]�͌epxޛ�Y������^�E���x�t�YZKl�j.#�20C���hH��']^HS1���{���7OPe�q'��rQԽj<���T$�[�N��2xo[�aSa��:����?��w�a"& ����-��̇���������7r��\�u����9�)�W�QI���+�uT�ڈ��e�cf�l"bŽ��d@wɘ�k�\ػ>UXU�n��Y��y��G-���^�z��E^�0����<EU�5�ވ���-���+��I�(.�@���z	Q��3(��Kr�]>a{s~ B�d��cC"C�$�1�x6�Ў����Jb�ߺj$L&��V9K�rE�d�r�)�RGL<�tt��ɻ�M����.��2`P�f��j����S)���@s�<��*��'B�q�f��xk8����$�1��g=���䝻"��m�z�ݲ��rH[ƈ�}�ra�lQ����M�DI��~;;)��z�ME��R�ZW_���Lj�S�'�_��Cg�H)����y%؉���M�~��$-�#���ep���8�*��"�D��L��x���"Ƃ��k��SE9Dޖy�p��tB�[�)���KT�"Æ+[2ر�k<�ҹ�L̛>���z�����^��dG�#��
w8�Oc��i4~�Gڥ?�uk�#������T;r�!=�9S:s����Ǔ'F���b��L�i�'Y��d�(����M��� ����r�3�
�^��Zv!� ��[{+���(�H��7�0�P�6+��g(B�VB3UV�͏�D���2��a���?�	�o4x����Z6�(l_�N��?G*Op�4<J-��]W�[zte�u��Ұ��q��<�%yjC�����`�:ؘ�^��`Ъ;~#�A��lM�ilFO-LŁ��.�H ��x������!֐㗹�@	��ZdsE�I6���d�G��9�I	I�~Ʒ�n��[�:���^��7�H�����m>��y��� ��^��/u�����2���~���ݘ�05�1�X�	�~��z�X������=��U�;�-���H�>}E����d��;�ZTݓ1��Մ~?v�a\�I�z��F�1^v��������+`k����[�2ʃ���e[q�S�)��Q�9>|TU]�I~�����>�\P e|W��'y)�j�ma�����r��/��F�1M�<O�Z�mޅ�y��Ld�k��*�&�]P"Ժn� �5��'[�G�^Z��Γ:��U��`b����%��:�����K�E���q���Zܨ��r �6�>�%�LX;�Lc"MVE��X�>�k�ep0"8ը��Q DWҋ���h6�9f�i.�bC�D��Gf� ,�Z�˖��=sn��+�"�_4��V��6��%{Q�P�c�z��֦I���o�chvb!��+���i;9ZP�E��| �/"��O[�m���s;�ћl��<|��+D���O1۹@p�. ����~z�u;��ǆ8�����Q1�@�pz���!5�m�z�&l.��4-�0�O��Y���G�-d�uM?TRېL84���5�J��tEb�dH�T����C�tN+iT߶��X�˴�<k,�I��:5�	��葄O����H�V��-s��ڱ�*����z{.'���38{~���׍�T!g�9��su��GUV©F����5M(}�uJt�g$�C�CB�8U�&���j{s�iHH���Cxg����x��ﳪ�N�
��My~��3� ��w,������5����WQ��D�9̸M��\��s'���<@�8����G��n�NSG�`Ǥ$��gH��i�s�@���>�)�D*lG��*���?l���/���@*|^�g=L!����?�2J�l(U�d�tF����
?��+��z�E��؉���`�h&0���FU��j�uU3
��~�y��j���Oe>���0<�����p��(y����4m�`�|AJ���e'��3Qr�n�Y�&<�x{~%2����B�1DO�j	�-,���+��BEV�M�M}��O9���q�D��/�)�u�$�~�0�mo�@X;����{,�!_��\^2T�~��H��B&^����F�^u��.�qO�m�q`�EZ1̍�̓��s�7\!��8z����s�ɶ��N��H�Ͻ*��f�Q�Si�)�F
>�jb���U��80�r+������ƥe�OB��d�kM��}�M�lZ�SO��aM�Rd���!z�K�	�W���w��2Į�����:t�"�{?5(�'�)��L	��g�<	\:�;T4v]��[�V<�#���3�-k%����񰑛S-ʬ�rRx��H��Y�s.\���|-��/�\�D�z��quOVU,�?��	�V	�����z��S��Q�Z���S�nN��y�-BΏ��Jɽ���1)z j����W���5ud�~�	�K�V]���%��v������JV��w��wh�sݿل&��s]@��<pl�'uo����؈����"q�۳�� �5�CFY��bY&�U�U=_�g��~��g��ԭ�܆|��:��ٻ����:��qO�c(u�$��~�Zu��g�(�K��A��R�P�D��N��+�H�G��4�aiuғ3\v� B��h�U�B^6��eN�'tV��$��h`-�eTcۉ�]aڒZ�inb�~Aw�j��,w�3����t�s&��sE��	$�#6�JM����������Fbeg�橝U�!�jo�L��<|��xUL��� A+�9Y������lq�/�i�>��6c���\�pIE��c̕^���w�	��N���5�eő�[�&��*ׯ�HF(=!N�Jg���_�5���ya�%�1-e��x���]lj�o�w���UO�|J<&Ҟ�I�m��KJ}��)a��K�`~E#܅�j%�r�q��- �湠N*3��uQ@i�W���m����>�ވxN\�H�.٧��ldg���2�x�]9P��r��k��f����a�&E��z~
L�k7�0����S��0�U�O$���|��'S���i+f���'h\��g�DePƔ��x��U>,i����䓤hO����3��^OT1�1����Uc�3V(�1~�*��������U��Tg+�a	�4. �f� 1�UW��,E��aU�q>|������z��I���`C����pFE|ʂ% Z�4F{آ���b_Y];j�p��\����1߁�Y\�#�8)
ݟb���H���8��L�o����NDQ��&j�F�3�F�Q����-f5n->}o��DQ��uk���:�8��d��T-4O���h@M���0i�6��JFĐ9,Cp�F�C�iIv�Yp]G�y�Lț�ƶ{xY�"�E�4r���`���}z������?��綧���<OK>Q	��Q��(Ipq�).�J����L:.� ���z{(ը���h�©�_���o���vG��P��4�*��<�;��_oM���t�ޭC_-rE�y�%%�ĩN��}J5Ɂ+QD���y4���!)闝� ���'&�1K�A��p���W���x�J����
<��6.�.���&��J�M��R�����Ύ�����3G	Ӳ���\�{}X�0��;�@Zf�2/�b��b��ax�����:���J[�eC�� �R��9D���De��f�!���
�1���V�t�,2���X�W���a��ߊ&���X)��N�GVC$4����y�X��B���J���69���i���������5�n�=���(�(I}���	�>I$��y[���&��aw���P.�����*h~֥�X8� ��@�m谥2�$m������=n]��_}hMd�+��J�0=mt0���.J��Ls��9+�E����#���VN�b9����r����őO�,��$�5\��I.� �"��m���Y|����@���6��3t���_RFwK��S�o'��e����pk�����ƒ۰&�V*K��JLq�D�_��?O� �լ��P���έT�܈���B�&1p�b�'w��5Hڒ�x{W��h�٢��78F5���ϐ�ai�X�Ά��,T}�&	���iU<�6V<.�o;�7fmX��7���p�L�:P�.�B���RV�^ˑ�:s���L�Q���,P��Ќ3n#a� ��z	�1���Rϣ[���N6�nx:�L��`M ��=���Sx�A������P�a^����L�N�rS�z�)�%�T��kNjL��23�2��ɑK�"�K��!S_�%#�!o8�_�1���|ۃi���`2�ϯ��
J�QJ~_P���t�V*35�nn�UE��H�ؿ�Tp��d0�$֡)��7�#�ޤ�ڷ��}�Y���m�x�珣�:�#S�h��qgPV_(��W�r�`�i9{'������a�b��ٿ���e����'FȪ�f��MHjJՎ!�`��`"��{69��lǈ�O5o�I	Lr�$W-~�
�	^�P�T�9>J�����fs�}K� �P���$tq�@�q`�����0��y��.�Eox������Vr0�ox�X���c��Y%�ߩ�����eau��
&�,2��J��&�����m3h�\�\�X7 ��j�pzV�����w����+>X�R�5qI��s�FC��	:�V�]���թ�J1���ͱ������J^=�NGmkT|�q�anۇ�[|������dΙ�i2�&�e�N�Yb;tnU鶚ÅG\��n*���q�@��jՏ�pܐ��q���q,1^��`O�٧H����$�8��M���@���`�o4Cמ���r���uڟl�`'����[�&u���W���,���Ǖ��+�,кʼsK4�>��#!o�����Pr�$�m���A�!r�?����	�"3
������JM��vPDgNT?��_'/>��Q��E�:?�%�8�-<��A���Q��}��7@!BT�4'[e�g�͔�κ.��d�J��N[���O���5����s勺�7�|o:=ϝ=�A�ze��|Y����}+�$��u��2+�n��&� G�Z�A�c#�Yk����-I}I�%�o�*C��� ��s	IS�"����I[iP0�%�t0-#pj�7�dm�
�n:�	�e��� ��r�]��{):�\,�RR�q��O׺	m{_���IH..��Xw�}��\l� ,lխ�?}}Ɨay"�h��R!�y�`V�n��9`5�f-1<�n/��{GYV��H���X���֨N�t	�2wgJ��RaDqHJ�G��O�Z��V2���&^ %��1��'��Z.�Tk���QU�7���;?_�c���cq�U��O�KN�U���I[�M0��-���H�����}����`s��.|���þ;ҵ�2�
'������ژ#�h��1*n����Xi�w<wWg"e����4$b���/{����{�z�/�=f�MQ��
p>���S4�y�G�%��;��y�=�U�������U[Jj�_w�%����{v���2��?��'�U5}�K��J¿-�\�<���fl�9꬝�u�+W���E/�\���:%�B@Z�����[�&��aqK��+�p�
1>0^�}9���5��!���sO�2�Dު<!V����m6(O�u��;����H�ج�����bܓק�쳖��߅�R�)�tp\��"Jb.4�������{g�<a!3Nyx�ΉZ���S��b�iO�S)a�:r�O��9��8o�%(ܰ�X�Kۃ��?���bw����mHf�����
�6���h���s�鄧�s�����R�� r�������$�������X��p�A'7#��N�T�D��|�"��e���B�M}�e,�B��/�5ĭ��E���S�O���ӂ�I��	�
:�8L'�O��`�����J�r��dWjJKK�d�>�,���7\�ZA�@�YaX�ڗL0.@#�DT�y'JL���$�_�b�5T=W���/s�ZW�R�~A7�Jm]>����}�~�2�r�av�cT`�χ�;sr��Z���Rwy8���6�^�JS��B��B���V�yf1T
[� ������>��1�nK���H�t��- �t�õ����&˪��Yhj����?t��[�ruU���״b�����њ����**{/��oKт�?b@*<�������������-�M�=���^�&�Pnݳ��nT��J������Vҏ0�>,SgҬ�JH̹�_���/���Eb�/7������)��)T�*%����2���V"�݇�F�o�Q�^�;s޶  ˜��n@�/�=�m�1bV߫E�q�S�$��ֽ��S��6J���R�>XD�VFV�6����c�J=�5�`U ~1<��6pB�3N7;��խBg?S���f1jk�'�֮
A�P~�OW�@$�A杦�ކ�����:�u��2�y'�|��(���I�sFu6sF��'�DAgd���褕��Q�c��p�.�*�BׂS����f9���nXw��A��^"}
�@:Z:�x��7S�����&_��*A@K�n���WҐ���{j^Y ��h��,m�ޙR6������qkSW�`G��C 1
�䌧��w-+{��c}U�B�������/#\K%�YU��૏�t�X@\rh����2�^_���4��3�ݨln���ͱ���k�#h�ۺprr閕�逘��G�cGD}�%y("�{�i?��y��HŅk�
M��	S���l>`��g�cv��v���
]w(:��!>T����#e]�h�a"�Z�d=�%��k�X�T��M���֢����6P��+"�d�hV2TX��(�
/�,x-�F�yw��n���ȫk�> ��Q��DHw��>?����M�h���2a�a�%�.0Q6	��Pl꨽�F�=5HL_I�W-M��I`�	�iW+k�]�k��U0z��+�ǙR��ҟ0�/?����T��F1�h��Ԍ�+���R�PG�G<O��W�����[�
�45��1��歋���Y��N7�n��w��]��	K�a�ϧ��V�������/N/,�_���;V�7�H���,h��i���ۣP*Us�n�U�t����r&rS���ʺ��`{��*Cl�����>��R!������ ���!tK�2δۭN8��T�k�8��
�e���r���j��Y�ץ������c�ܢ���1�T��z���K!]/׀>xs�h"� �"R����/\9��x��3�.p��󶉅�X	P�`��85$!����4&Mݱ*����5W�%J�NƢ�tu8����#��}]�鷎�B�A�R�	����>��b���=���9������R���o�����Y`�D�W��%T
�P�1��R<|;��?�6�-�gʃI����1��j`ϭb��9���x['����I���P�:`��%�`���,J�ٌ
AK���l|W�a����U��)I\@�BS��y�g�3pK"��Ɛo#zVg�jڅ�S�/����h��,�ia ?���i|�EC���m��L��,L�,�o]�f��,��q�]�Y�-��w�_��kH&���eλ�\M��V�N� .V�i� ���s��룽��2|��Z����⳴�7K���~K9i*f���_�.{73v]����h�H��c�{��HFe�{�'>��2>�s3g)�����W9�S�#R���PX:s��e�Ӹ)��B$ǃ��2JF-��O����Y4}O�?[��F}����{:z5�q8�0�_}DG�nk(��LpGC%qix��()�r����F�O�#О��^s.n��I�f��^��(@�:-"4��Z���ZlL���@��6ǯ���#��v+3����z�D$M_7Ʌ�g�ذ��1��F1��-{Zr9�D4���sP�L�K#���g���ךJr��c�~�+�G��Bo���^����[9���Ӎ��f-���Q�h����qf�k�ϾTʿ�8ms7�{g�D���V����o���E�����U�	��=i�ƨ
��AwG������;yP}�0����( ,�
�t�c��O��m �l��2P�h%�2�O��wK��:V=X-ݗ�W:R���-Z�yķ��� W%e�b��\�>-i�q֙��l�����vK��F����h.kST�׹�V�#yU��k"��m��*=KDл�j����P
]��9�C��o��3�;m|�R<Q�v�x�Q{����ʁ�y��R�Ff�N+�@;�R YK䜬\&UGb8	��cž��0EBmP��l0��H0�@�Q���1���K����p�Ռ�l7���5=��,RBP 9��څjO��W g�D���Mس�^	{�����/1 n�Z�Վ�Ko�9�m^��i��j�q�[]�"a��y����W��/}S;+�k��FR��A��S�d,�Z�z������w�Nyc�	,�9:�B6&������)��>�y�xj�`w�
� ���H��i�R�1���7�PL������E�8�@�����} +�9��6�FҨ�)��cn�S��U�g��6�	-q{O�i�Ħ�j��\���/d��\[ị�j���.|7H�k�
G~R�0�<�bR�=f�x�{}�h0"��$3�\wpi�&���Z�����o��]�C�F�~1�x*ѷ}�[���?��q�nRgc�6�[� \�e�\<���t�}N�k����C]��W�`^�5�Y�"J+�&n�o��f�7�n��A�}�5^`�(×AP�]�R�Ù*��N�z�]�|'d��@[�W� �^����>xq��=E�p8�EJms.Z���@����s�G?՘|�
1�R�dQ㏛��!n�鈄��̘��t ��2����@ɽa������L�c�{��.����:N����qkP��x:Ͻi,s�2�jhu�&�(ɉeS�8s���x��X4b��h�-,Y�U���>쨫��n2k��H�ۨ�n��Jqdn�\�~��|�w�{�3|ǝ��I]I���4	���<#o#5uH�Tz-��� ��1��h�m�߼�qᜓ���V�#�nVM��fg�VqM����s�!���IE;��)�«����W�f�>TF��޶WĄ�붊`�-U��<�H���PvN>�e���J8j�ʦ�o�D0��UO+?�7������;�����({�ϓS�,���9���CZ3�a�E��Sccn�C��#�թç�,���+�&��&#q��Up�Rʺ�a@���R�� l�J��ޚҸc ���������VUX��A.������cq
�"9{p�� ��c��Z����h��t��[����gu׫��`�S�V��K���Y����5�?"Q]��㺷�@�ק�}nwA`7�����鴘���@�m���{��>Wէ(�kf(�?�1�S�&Y||3{�U�N����@�S���~�������5AE6�ӿsU�A-{#�(![1�ޞLr������H��7'd1�ۑ?Lgl��eћ4~sY'h���8K��kJC�*&�f╺�Ui�E�C����d~=���S.'�Z�<����L/�"���y�]�i�+`�Jbv�2�1�<?J��p2��ܸ�@c��$Gq\o��.�c����J�z��]����]���E<ܲa���d9'�L�*��%�e���lu��@�aT�|�u-^H��Tn��Y-�,ݡ�6 �ag�MRX��7g���y��	��,Wn�TN���l*1�Cp��_��@ޒ���g�۫E�N������Wn�-��)%%�W�f3[s���"W�o�s��]��|Α��v��z蔏��"�����ὠ�,?����׺p@{Gr&��$�,�Pc�K|3�?��(��� �T���S� �s\�k�;�z��r#1��X�����X���\$�Z��]���T���];��z��o+� �b�v���,��}�	�]���p�2�%RS�\"H�6��%�0�������C�����l﯃�d!YB� �a�ܚH�xO!��2�rl��
	H�Sލ�ꁬד��W�UF`��Ew�j���V�RթX��a���]�ٽ�O���ie�5aꦃ����i�:��U#YA����K�|�d&�h�T�hF��mu��}d8Y��0��m��)\�"S�>)1f������Աh\�п����qFn+�!��&�_� X��	���j�}�%U�1�i�>�T��rѶ��m�rc&�!#{Ո�J�!L�'����lf	A��|F<��r?k6���SW�Ȝ�so�ݞ�;���@"c}w�˗C	��3A�)V��a;8���p�F�J����z�$>�V�~F�նK�U����_��عZ�d������������jq=7(��@A���y��PœW�ˣ�ׄ��"�UH��c�~iq�(5I�n�#��uWBr#�-5�}��0i@G�?5�
lǍ[�t ߢC.�U����8S��nU\���$1�븋�_ 7p=��`�;��c��#�0}��M`����Z��ϳ�qvR�1�P"�P�F'Du5F�T4�����DWܕ�Bn�p�� �JĦI�v(���t��w�b�j�n=̨pY{'��&p�2�hmڑ:b�\�!!)c�h=^�POC�$��L3�r�]��*��<���d,7���z�ɪf��̇u�k�ll?a��'�]�?wF� �$���_��1C�YA�/����w'YN��J��½�&����'<�Ѷ�b�	�)P�W �*>n�%�CNł�Z@OE� ��䟉�z�&�\@�_|
�˨c��yԖ�֬��$;y��Aj�7���e��dNq啠~�]sH[��et�6;�SR���-��q�1 ��{���l	�,�ݑ/�xK'0�Mt�VKK�������Gk�W. ������_��A�a�mIUv���Xvw��Ϥ�H?���ҁ��z��&���q�H��V�>��j������k�|�bי;n�` ��Na����qM�I���������ĒT;IH��1�f�-�����\�n��i��c���=�N�/��L�@ݶ�����{�QT����F�z�l�ָ�8��Z2zb�hc,���WD��$���RE��xm��I�C���F�|zC�f��&[8;�IoC!M��	wOg��i���2<�mP ��w���t��e���Q��ع0�N�Į9a2�CL�99,���V����}H���^��!��'Z$8�U���&&��B�`�f"p
�>d��X*�P+cŦ�5	��$4vjopw��gB�ݦF�ZW�au9Up(�,�����e*>�>�aH��:�v�s�@-��)٢�i�ah{P��zd`��~Ɣ�7@�S���Q�+a�+L]?�v5�G\��0��8�C/�p�:X\9R��E�۲�ձ�0��h�G���CC�a�8x_���L�������Ou4||e�r���b�q&�|/&`�
,�_hd7�(�2֞�[�|\�%@a�P���:�,��*r:f�t�-P^��.�$:�k���7�xl��;\'�g�]��yM�r^��w��X?���z����dc&�zy�HM�N��� �*wy��umGh'�:�gB�D?Q��U'�h��V�@��e)�,�n���;�F��K5nM�ڜ-��ʊ��z���꒖>�*�X�U9bg0�z��}B�ġK%=����/+/8Z�j�?B�v�4�����7��R�8�S:��m�:�/occL������Jkb�������[���ElXUS
�����O��_�kiM�����3D�~޶$]'��.��[�h��U��e��
�^�����>%lp�nF��p	ƻf4_L6>��B@������B"<�>q��g���mK��6x,���%��&�3��dl������s��[� 8#���Q���&��C�D�;�7T�<R�Lf����?��B}�!�uc��2E�A�R��<C�i�f�$oɇv�h ���K�R����dA�Y63̤�����U���Nd,:v�����8��D]h����!Eӹc����-��	U˙V��|�u�z�pި��p��g��Wh�	�0����@����,����g�+�t)�T���T�W�ka\���+7��K��E��m��)��_�o�O(�᥿�A�:�m)?��^@�c�S�.�q@��������_P�v��y�L��(�?j�NsUA�m>�d����0!��G%+�&���x�0�7a�6�Ut�7�_qB��e������^�g�஡ܭ|EJY����-�BAl{W(�nA����TPP���V��o�*]Y>�3�����������g�T��2MI1���X����E���J.�2"E�X���N��Q޽R_��4�G'�ҳ���Iy�-����$�5�QMR=��r�z���W���쬼����G2!��	)�X�Ƕ�����ףA����@�1	�I��bt�=@�iI�>�W �%��iOqs'�1&G�V���]��:JЯ[C��~~���<08!@cE�V���H�n��T�-��EE.�A��<���gu8#�z�5	��6��v�\��
O꣉'j6��S!9s�)v�,���1�� 7�/��˚�$3Y�/}yM�ҼZ�-(<K�1}ġ�^�λD�[�Kt���>k��@�|}��kfS�T$񍘻��>�i��JZ�JV��|jf��������=Q�ob��h�ZS��m�-�[�5�A�IDғ�#q�O�2����Y����|$��8LQ�o�@~�_y��x%���}��$'<���3dQ��u�8����ޣ*��i�p�덇$��i����\�Q�bxG\m2uE<OH���s�X�䝺�:�/����N���ـ#��k�6}�!�<��3z�@{�K�M�A"`�PE!�H���|�ހ����2u������װ��ި���W��I?��U�ҥ��@��m�;��{�~�:q�PL��#�@�9Ӥ(.�����i���J`��L�@Dv���oY�t�N��)�?�&�m�c �\J ����ZA?jp<�O]���Ts�]e'w��mG'8��6�����譞)W�	�UJ�O��wu�V�$�ÅZ��b�I�����Z������(�w�~Peb� h��J}�9�}�2^��}�Y.� x�>����l���v�'zۃt���)�gD~o@+.G�;Y�H��9����M/�Z
,_��U��Ii>�*��,��C��+l����8lu��,7��*`yX]LaM�
��%��ȉ�0O~�Y���� ��e�����T��>�b^��])���x4p���1����vy���>$�����%y�s���S�D�>�':�p��׵ʈJ?Ҝ�A�#�#q8HNe�|	-�n-�J�;�� ��������M|�&�T�E�5 tCe���	6Z
��g��iʟ1<���9��3X'��Kt|z��0~<%r��t%I��JB6�ɢ/2�k���H^����A�����j w��.�۷�G�2�zp��c��+�ۉe��ei?�uZ�}l���n���+]�3�a۹C�tZ�
hJ-��Zi�+ۋ��e`C{�.��T���!�ao���w�6B��"l��YF��Y>��ao>R��߻o��i�����C���7Źq� ;)-�{΂&���S���]�����^����B2}�-�#�:,���w{������^C�����*:��9p~��oHDw��� �ɟ�$u�����#ͼ���@A�0��ט9Y�'��f"��~�1O�*i�Q\����2��9��D�L�����2\�u�&=��Nꃇ�"�d�u^���d
�j���R��T�cR����n"Y�V �et�����ٿ�ϯ�����;��%W��b(ݭ�#�M+ ������>"��#'�7v6轋�v9�#&�s���t�9�ttk	2���6BG�q�o9���������Ԕ��^�9��>�R��I{����*:B,ٴ�g��9�#$7���A��=c��U�@:��%�ߩJ9����I�x�Y�<oZ�{�"dA���	)H���a�״��n���`�>g$�%;�Z}18s����=@��],|��Ɂ�#��� u��x��@�6�za��S+�x]&��"�[4㠮��*4~���mź��M���|���A��IX7�.z^����IB��h�)^y������L������й/�y#�vf���`���ޞ>m��a5�O{�"��[�M�0���_�_poA	��*ڬ����XU[3U�Klzɗ��O�A����HMpQ�j�-}��p��D�
��Fr�⥑��>�fޅĞ(��-Z׼��ve����6_E�[����4����(��m*OE�/����l�~���@.�_�(��j��f �2��s�>��q�;G.�,g���6!��
�|M�w{��.����{��O/-4��^:�1��^�ί�n�����[� V!��w��Bt��#X���5��+�T�t�L��/�c6W��e^&	Bj:���	:Bֶ�[$9�o��D�C�������ˢZY�����SA�Sm�&,#Biǡ?�k�l̪��qC��?R��J�!_:��Q��'�R�v?:��wi]L�Q#y����̐�(6��?!�
i@p]%
 �͞l��d98�/X�PI��e�ų�^�FE�۳�C�x��`�5�W�{�$0�b f����{�=�'x^�ym���`��M�J��ڑ�w�.ۑD1)Vߢ=gcG'��ry�݅��ql�X�?�E��D�@�V�c	����S� �'�f�P�If�A� �F%�����e�p07:�^����q\m)����Mٿ�\���J��I�M�=�C����P(���+�3SI�*��=)u��+�K2Ѫ�{᡾M�z�s��f8�;.ӏ~E$�/�u:��*C��<��0�Ӈ��4�>�f�1�X�!V�%X2�d�75��R��入 �d�:��ٿ �B�3D0Ȋ;�����[d��
�7�<�0<��vg;�(����+������G���!�h�4Xr9�o-�x9T��q�d�/�0�J5p�����ۀ�bWN�J���x�ۨ�L���c�D�60���Ѐ�A�����3k쑴������[][n�E�d����f��v!���!�x���v��uw�]��LG0rР������$'C����
+��~�be�e��`��T�h8��yLGz{�5��WI�	Q�;��C\�%��W�>m!�����@*3�ϙ��TӖ")�q��hiaB8�Tp�ڭ�@�g�`�į�Z�J�דi�'���Y�oٵUG���WDc��H�6`�m/""dl���	ˁ�����CS�G>��L��W�_9�W�+LBtxB�����49r��̬di�����|��"|��_����N�D�O�;F"Qћ�x�j�.�<f\���P�p�=��_❷^ژ�X}9,|i�q$�[M�:EQg纯��{�̓������}S6��q�)�q�i,��LX#h�U����$^L�ܟg���j=}��x���T���Ux��,�
ڜm��.;'�Px�r-����J��q]�/Ie ]Tj�K�v7�?FK��d�������ɍ[o�U�c�w������%�T�)��<�����$iʓC�#�yfûϕx����^�=����ӳhL|0��J�t9�]m�!H���_7���^�!�S2���ţ�K�f~f顊�J���x[?�\�[o�<�1؀�ת�^�G~in`^�O	-u��0�
!	��
�(���W`G����G� C�\o-�0����-���^���(�I�c��4S��:�e��:��f�������`W��(G��[ϖ�Ft��0�O�R|��~��j�	*u�W�\I/� -��a�6L �"˰��-
d��|��&��C�"ѽ���UbA����t�Y�����!���٤�*�����}/΁I}A�� ^�Ut!@Ng�?�i.��6@^�Z���:�;W�[pv�	�{�n������uWҜ_��?��2=�fRbv-at�c�xTpe*�]@�5������i? ��Xŧ��]��~��X%Ϭ��X�ʣt���nr�*b���j�g|*D�(��NCM-���7��/_�k���=�S�Aq�7ܛ=�,�J��S��I�?~"0m�6��Tm�9�q5�UV�I����[==�?��8f0]Ȫ���� �$���,�@��RA�J�O=Nb��"��UﵘK�.�5Σ"��T��X��4��	����[BT"���nk�^o���]�:q��\�yZ��%��D�,���������4���ʷ"Nc��4���aԔ��$��%�V�^z�Ά�w�|�
��UZ`��X
:7z��i����C "�aO��&�%�9!S\P��,��ȟC -f٤x��dPm�Pm����{�x��$�В
��ߨ���)��9p�n�D�(���M�Qg�HY�l�#� U~aND,�~?��XL�Rv_��,MS4���q�E�Z�7qa��L=�Ea�Z��˃�-y�W��T�������>:����@>@�7t��.�S�)�mQc���)y��������fD�|+��'�ԁٸ�E�U�C���Qe�Pj|�B��Mj��wL<"l�����X�7Zy��*��y0c.�U9��@ �g3f�<Y�n�I�>~坸�u�u'
�f�Mv��+�'6S���y8�g��n���u7��1�����14|�����p�qs����o@��(�HR��X0E��N8G�;ކ���L¿C-J=f�1�����B���10�AsZ���Z�9w6Ta��JG��8 �_��J܃�2�[W�p��%��8a$��_�����\�D]np�H:�c_G�����:��p�>��(��}�Pe�P��@m|�Ǝ�ڽ�i�+i,�?ǒ�L��g��-�'g}�{��H��Qn_/k>����&�b�r�� �5�3�B��a�6�ο*yE��ב���T<������r�O����콼~SUH������`����/���Q�*g�WW�e�i�+۴ �
�JD�����O���u,��9�|�x�BxbfG&��;o�f�d3��<��TZ"�-;��g�:�nO��g�~
  ���: �����q;�~���h;�q~�A�r�!�\@_N;�h��Վ^fN������/Yva?����������X�w[~�k˄���ݍ�#Q'qzI�Ґab2�k"0��iϦED�> '�ïMG�1����9��o䅀�V�q}�: ��7��M�����1eo�u�u�NMCM��&������iU>�Ρ��j���{�cg0�F��3��m(�^�4�vy��O`i��V5Q�Eet������)�, �;��E�JZ�.O��k��݊�
s�.;2��m`��|�o;t��gI��vUp�t_ ��'1�.;儸[���Tt�Q~����'����K
�f�!��ß��|�� y=Q�#C�9��8�p'%䍪$�,`��R7���2�`>��w�o�X����<�g �Q���� ��$Y���;�E65��&i:dw���>$ec�R�T-��:��������)���g>ų{�0���C,�mV��� ݘ�)�  �#S�)V��wԆ���i�w�#��b;�g��]C�@#��W.L�D��7�9�\6P��������v��D�{k�*��-�	U���gD��o�Q+��rA�j�A���WI\�[���΢9��ز[�������y�d�=v�0����)�s�����I�C�[�G�ÈM�ŚV�c3aqY��D�z�!�vG�q勛�8�:�3�7�Ra�<,_����&�SZ����(�A��؃I\~��h� e�!�Y��;� ���]X_K/F�цơ�;��=���#K<Y�X[�O|��Q���ģ'�+�:�׸�ʵ̥����v�a�}٪2��íu՟��Ͱ��{r�9S�Y?�W�I$e��bXC���)����E�ȇh�����Hw' �|���nC�V�'��[��Nz����=�سv�J�0��'�s�
s���>e�UM�ǜ�������e�"�>\ǥ�UYZ�^Oe�^��}�o��Q,W����O
Fb9�bՅW�Sݮ'Kը�Gi*_F,e�lm�ԚF��ֲq���hc���x����0s�KFL�D�h���H�Rw���~ܬƿ/���!���_Ԍm��y1�Y��=�~���ـ��n�p�?��5kN�y�'�no$��x{!���
�ňR�j��z��u��to�NΏ{M[h��u�l(�ú'鿎2nU��D:w�6��dш[U�2n��;?U����{t/H���/�I/*��>��S����j��}~wvzK��t�\��g��[�<S�����ϵ�W��*��� �)��<e�j
�g���,��@HK��Si��'����m�fI縟i���4m��ٽ�RS$bL��򹭬'��c�W����1���s�X(T�������_��	��rrqd�Fr`�7�`�oZn&�G"NE�iFC�d>Z,S���A��X��e���C,���NEThj�'#0�WL ��x��L/��f�8m*�@�4rR�	���)|��S���@�E�\b����~/��C
�~��Uq�$���d[���1=U2xdj	�`�֪|�MuUPSahSQ#l8�j��yö�C���S��qV�(,&���Е6P�?Yo��f�%32y� WC y�G�m��	4)�$���$�}�8��{�;���҉⃸|w�)C<�tн��_�ۏo0�i��A߃�FT��G�#�!��v$�_,�	)7.M�iiٿ�d(r�� �B��}�����Z�Lz�AP�^&Q��$��}�=���m��_@ᅃl��z�����u�\��h|,Gh���D��i�Y��@*�q��4��(F=�^a���X�]��,�\{{��� ��s���D X$��!:���n�=�4�pcY(~���z�3ٚe�B��vI�f�׆I��q���]��\{9�A�� �ri��_�c��-�y�4�N2���D����������Yu��'�X/V6�edE�1)1Q��7���
~�A�}6��"���أ�dC�p���������T�B�gL2@g-=�+3}��^����@A s����ֹ��p<u܈zM�[� P�nd��\q��DQ8��-�p�����C�꺄Є����`�pX�P<ŦF���1w}s�!}����ԻL�dݣp���J���p5.���pxM�Ř��W��J�i������ҧ,�i����t^D|�!_}tu}`޵	G9ǉ��9}7��lmv�X�:/8R���
�ÿV�a���ˋc]ڪ���-��UJ]r(����CJ�:ﮏ�`�V<
mN�J1��.��i e�A-v<��}6���\��H�L����p筏ܘۦ�LZ���V�[�R4$?	�0�d�
��tC��FjC6Uf�;_�>������&�tR���ep=��	� ���x�n\��D3�����^S;$ꄪޢs. �[�דҠ��b�4�cH}��ߙ��.p*��Yu$ڦ턄�^
E��9],�6�o�C�;uh��ɭ�5ѱI�����B���r8-*��a8/@Qa�L��z�l�W�FG����=qř��E!N����L���蚪��wr +b�)Q��{j���O�q\<o�wC@�����kKqgF�ޜ��	EY��k���x���4�7����W���n��`ؼ+<��`9�rYb滴IF������%�C�M����3#N��L�kB�p�Yt܇P�����%i�@̄wb^���� ������?���Ѡܤָˢ�4�t��w����<�?k��Y��ޅV�٦x�F��S�V����&�)��:�F��\��y�ٓ�]��So�$�P�* ��x��aG��:
Xs����*�p���F�c���5��)�/��8ᑵ�lbv�	�]���Ǫ��U�Jٯ���ca݁>���ШR�St����������������������w�9)�_x�VA����6A������Q[L.���R[^z�����s��{^�6~V�MbRa�J�,,Q.��?����h��p���14�O�h�����9�.�*�E�aVrY�3L�7���G�7��G��;���虀�n>�1��{�	%xΈ��2#�Uye��%�!����Sj���/}�jx3�UM��¥��ׁ;U,x�lg�~�_�!�\���$�/Y�yc|�^WE2�b#J�|���hWE������|��Fjsi����Z#~T=/�;�v��L0�*�������K�
��}Y>�}��C�P��l�)t���9���K�4�s֕��^���
�! ��� ȁ]�����Vq=�m_���`�����͙nu++F6I�?u���W�Ih���|5�9$�����sO�X�q��;���F^�w��Trg��P �)X}Y������;�'t���4%�7<�#�9��J�h?E���9o��eK�
'e��OXYbBA���1S�����\e"��j��.-*y�;�N(��'��o��%(গћa �-��@,?��⠔�a蓇?�(�Z$߁��_���U�9't����*���#P!�V��&����,!���)ހ��W��j�{J����hGf,��(���n�G�Pm��-\B�o�e'Ȫص
�_"����r}!�~���U-�G5Ѯ��T{;qo뚎:����P���u��S����^��&��a�7�Jᬝ�<�	�� �=�u|pi�e:��lt�J���Z�2���j�^���� �B���{��e|��1R׾�+�g�b������%�g��%���T2=p��]Ґܦ~1�*�n�W8�0~�CǺe���ۦ�ed+�ӸI�	'�����nx,m�-{q��VË0��@���)F�jc?�tH<�S�F��L���u��R�!��c!x����C���攏���@>�Ň���~�!�����O���zӘ���0�>�T��C�*�	�i�/���^���ա=	s);ZVù�*�@a��v)g�H�֒��g
�9t"|W�'a��������t���4��u� �҂��:�|��J�4�+ �2sN��ظ�����{�Ɋ/��]�AD�����4<�z�������<៙JM|ن)� �#2>�K�
�9�3�}H�|����a��]_�E��[�>u\�]*7� ��7�T�6B�v�x}��A� �A��]XI^\z�RC�W�:����(= �@4:�.�:+���D���\ҥ����-��VbںObZE��0ub5�e�"	�UC��7��3:Y���7z��y"��ק2��ڐ���6\�}1��?D?jz���
"���K�H��9�_u���sN�L��U���}$���ha�40�HZ#
����I���:���R>��dh�ݳK�㏕ߝ���P.	%p��z~o@��qx�\7��xW�<x�+��Y��r':��HTz�~��Yv<r;D��ۧ'��8�5� Gz�� �B(������%a�\ʿy� .瞰��GA��r0]�`���i0'{X�>�rN�x�����~���a���9�%��<����F��R�ZE_���	�� B�R$�1�%&��w`(���+�B����6�zTSx|���44��%�ZѳIޑMT�hK�ǉ�Q�1�<��z2_���5�ͽ�oqo��4v����c�������]'�D�xWa���D�;v�Lv�ˊ��XuIX� ����}=<k[�����$�L�7��X�mؿ��9˃���7}��q�hBj�eA �Ӎݭ��vUgX�k�d�=����KV�O2ԇ֠��.�5���ih�<R��^�