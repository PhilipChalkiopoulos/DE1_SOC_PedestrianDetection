��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�kqDL��x������Td����|�{k�#i��H��/�d��-B>
o��t,gb���M������Bd`���Z�c�Y��N��\��$ڧ6,Ƞ�����H���Ѳ]Z�X��v���GqW;r�E��s�+{B?��,��ܯ����ˉf��2���Y���ea孕��"���QF�Gs9l�M�);�k&�
6����.�C+�lC�h�����|�6-q��k��f���0Ĉ�u�xN+7�/�����׏��)B�}��u}���xU�󁓤���՚*�I��8$����pɖ�xE��YO��9�Qv�E�H�ў��oh�u\ɜ��M�<^u�c�K�Q�����ڪ�P�C��	����0]��dU�dΏ(2;ɽ�,Ae|Z�>�ZYЬ/���:spuY��cY?a��_��dS�)��0����@�ݢw�w"|��� Ҍ_ƒ��JE~�M�`��ZЮ��.3��h��m�+��Ĳo/+���J�sϙT���~�1n�w��5��LQ�ŇTv�~/�[�;� �q����V�{C]r���D��A,\g[+���'�YO�ꋼ�Sd��;��2?+�:�RT1�]E�>-.�X���"��ʵF.�N�$�s�r`B}'�%9F�*b��׋��!�Q���l�Y�q������uӉ_ɉe�"�^��l�IA��~f�x6j2�.�k���_�)��zJ)�Z�hE	9�Y��;�p�w��Bz��J}�#sa` �mX�/�4 ���j�$~r���FD�ۡ��4�f���- �3�B#���8�d'����(2��v���m����Ӑ�KQ��᥮�:EF�*�}���Ό�'�3h�	��,���(��-�x�v��&�c�@�J1	�9o�g�g�*\���F}�B:�3CO�ڬ�,׈+��EOi���yE��Z�_6����!RP����O�J/'s�E< �f���MD��m����ch����7����{�ꄇ�ԯOm�M����
��J~jZ��K�L_/�ε�B�T�Mc2G.Z��k�%�/��?/�H�;}n����4�sS�t�kv1��<gUq �P�x�-��eJ��ȫ$`��dx�~Xd[Y��,Gq)�H�dx�r��Qۼ���g�B��9tg����VtM25�p�9[���A�@8�h���&�e�,�+�ɫ������.�'��!���-.ټ�H�:N��r�#��Y#+g���C� xi�a=u�� �Q-F�r��j�P���/��S�@���Z,�t�H��Ȩ��)�'��$}�?�J\� ��bu�ݯ�����딭�5��E���X�Q��$,���Kf&7�ӿv�[vH*q�",mJ�H;hծ���}�ˆx�\��p"���ħ��r��3�Ww��ji�������������A���|��q\(֌���ˆ�e�ˋϖ��x��T�)�(̟痤�U�rg���d�;?�^[��T4a�6\�e|A����0�D�+�&8lyF��:��*g�Y�vt�ȨH7�����Q3+rD<%J�+�1w~nq�l��4^�9G\?�D3��a9�s� �u����<0l�WI~g�iQ���p�*4M��q�������	1)vV��y�G!��6��aA�X�f,�������|& ��X�� ��Z�ˉ[�2�M-����j�J�W����(�u�.��zK��N�?(
��u�P��	������X�/��?G��A*�ݓ����(��&��������ϾQm󸄠���E֜B����F>���q}A�O��;�(�Ш�}��<�wncؐ�~�D�o�n*��9�3ul���h1��}��w��?BE	�~�ܧ�̆m5�	�ݗ��u����@����N�ؠ��ƨЉA��<[G�4�Ref)w�CD����Ye��(������g@�z@A�&�a�8r.�=oc~6�R@
;2��]��d�%�a��7k���h+!|5����o�I����7�E|���s(dy����2�����q�.� {��BP�ң��Vf��4�p�߄����1��?�E�T'W�W�ؔ��tg>�}H^���V��@�J��N��;����)٣�d��<B���9��T�$�{U2�4�y�1� �9�lM�1�U�#Li���E.8^��a�o?�<�x�)
iwi�G4���[N��X�e@����u��	���cC�>���B'(M���AC�pi�V��JNgx ���q�������v��ͫ���)���4d4}�؆�����p4��,��Y��7�&�Sq��9��YH©i9;�.��|P�q���j�糟q�ƕĶ�3����8����bgw�h&���E��*(����K�-�E�E�E�WMqI�~W�)U�܂��ޠ����]����m6CE&�9J����Yp�H�> Ow��:�"wa�-��\�iWS�k���� �J �]�-�u���<�
<��N�KS�3��A���tx���b������&#�;�׼�q�����ՠ�4�W�i��`�qZnV���xdD�)������B�o����n_Xز���1�-!�l�F��b��)��F+n���� ���Z�/U��OE��/�ɼ�O�<7M�V�z��y^�Hrk�t�a��m�pe����ju���S��I�&{��6�k\�.��
�o���5v���{�x@�� �<&�M�
!9���T�uU3lk���;�T]��zS��2BAbgG2�/�?5��ˉ�I�ݞ5ێ�����ո�dh׃�."���F+:Ӹ��f�a��FLZ�ph�Zȧ�������e��)C���G"�1�	����2�̗̌�✜�9��b%��:@�����\`B����O��&�9ՙק�j���b��0���o=@��ɌR*�&;��ߢ����V���o'���D\$�ݤ}��5�����Z�^����@��Q�h�s�-�+:��S�9��� \y�I�*.pS캿�O���i.v���Y�.X?	�4���xxټʬ���s���6��o%������eݟ�Nf�$�fyC`�L5},�L4�34����CC�&R�$
�J(�y��y!BM�h��{����ք����J���� ��a�Bc?[�B���Ѿ�8ṕ[�:>�*��{#i|Z�RL����Z*bo�z�/�5ö���w���#��oU_.�c��p�٪Iv�AA��,aY�����X[���v����T�cމS�	�i���em��='��>Ai�����-�;*v�w���������,��φz�`��s���.>�Ǧ==���;k�'/>�(��si�,i���#��>����A}W���v��(Q��@@xᖺ����1J3c���P��|?�1��l�֐�F����Ѩc^�O�='M��s�=F�r1<3i��@��Ɓ#�Ɠ;�d�,�EO��K5[V53�
]��r��Vk��o?����^�co�X��x���f�n��:<<�1R�[���{�4�<B�5Os[�RѴnЄ$���!��,s����)3�0W�̠�x?�����ق3n+�*�*r������:�����Z5u�[O��_;6ҍZ�[`J8�����R��N�\��SUC���4�"$utZ�tO��)'+r@��$��@�3Z��򧙾�u���84e�)nxz KX>Č���]5U`����&���#��s!����>
!�j��"œ�Qx����h�M�s>ǳ3͐�d��d�ĒW!�B�� ��s̎V�`���g�g)��TLh�L�P:�����f�`	��&л{�l����X�o���C��2l�U<Γ�W�@'_1��m>��֐�����!�77���̠Dͫ�F�n4?v�M�b� ��pc3��_2	75�"���~8������?@�R��68�c 9�bP�׵[�A�|�N��E�pA�>I���Ж�)�0�������;k��L�$|�f�Vy�>�����#yR��l}��D���o��#J'J��*
H^f�hC@=�w�H�{����L|��p�c��|sD<��C�.��e��q�C���^dQ��6�,��B����Ws���2�b��n�J{l#|�� 	�cK�����{�<�4�p$�� ۓ2�F8v����Y��R�
D?Q���׼F����9]�b9S�>���l�-�����n
��}6����Y�&Me�>�D���B#���!�?bly�W#�b�V���	 rb�aK�a���
h���9Ԝ�K�`�X��Y�e�S
^��[�5O�"z�\��n��=�2.�\1�zW�x]<��"�ş�J%}�D�6B�q'ڭ��XD`�_�P��G^πOt�cy�>B|��Pa��E#�4��������D����2�jS6��5���U3���0J�ד�l�<!,N�� Q*�1B�F�c���P6�#5Q6�Pg�VE�l�)��S26Б-�`� �ٓ}}�˪���Dh7�u�<ܦ�Q=-�<�w��p��Y�95֩
�����F���t�2�̄P�B��x��[qt�j����+���Z3��%k`�ۛqw�Џ�ƶ��U��r~��:^�����u?&)|抵v�g?��B�MVzb+ŉI���Lz�{��ؚz����͗�v�l�|Yv���(�����?�<�ٱ�����~�x�Py[\婼�3�Y��*���u�د_D�Em���=�FT�ب=��S!���T�?(�`Ix�M���V^�p<�c���ʟS��~�|�Ľg�r�|�����)���?=�����"���f86��1�/��N	��8�(u��|����o�:���nW�0j��{(�������\])Py(�H$�&6qN�� gj*	U
i*�Pp�S�'{-L�
1�_S_�8d�60p���/R� _$����zx�/W$�qS!�:ْ�>�{��/u�z�
:����Kɏ>��?G��;��*κ��ˎ=s���TIVT	TCJ�/�ʛȰ�b4l��nm!�ZG/���>�3�a@�R,�������՗�iUV���p�2j^ �E*c\+�Xܘh�|�ILc1�6��L��v|���V�[c�`��ʂ���ݪ�C�$u}����ؒ�M��&�Nc�LA�׃�9Yu܁hxj����@���.ϩDr�6����K R���>���g�O�%�������1���Ky����^��<38ۤ"=[l���h+b]��5,u�����y!�֝�7�ᱹe���MD��q��GPM� �[=,�E�Bl��UpD���s�V~V#����M�@���hݓu ��x��Z��ċ��y�8r23�c��s�i̎F#��=���|R��f �֔~w�hpkҡ��t��C�������#��.��A���ܼ'�@]�5���0��N9�G`��
(&X���ENK� ���gժN
��2$?�pd]+@�Ï��Ͱ`!�_lG�Q�S��Z0�m	±a�Wv���x�Y��E�����N�������wF�C�z뢈�t����?��|��$��v6�U� RI 7K?C�dAi�D���
112\�m��`Yi(��Ԙr��?V�f����z�)�h'�� ��ըU��Y��"�N8/g{�d&Vau�4R�~4�:N��,o�)�rtO�QV�\Z��Oi�~1��ݼ"2���C�ǆ5�4x=.��ұA�&cH~0b6�fwVӃ�nV�H)���Y��?��;q��� ��CAU<����F�����7 P�T�՞p��, �t"�Dr|a�c�������72�|��bfR*E4�Dn�|^:'�/�a2�� �.�&���ڗԙ�'�;�Y�d���~=�rD�٨qd8lYG��S�����a����/�������en��YdxqCڤ��r��3(����V���-E;hC�r~�PφTɃl�3�Kj*_��Ҟc�Z�06���AH��MC\9�z�����=S"�쿃�O$=�Xڐ���,5r�Jy<��t'�G��P){`���5������hVz]Q|sȋ�#+��>A��ˀ��vGCFPY1Ľ��L�(����Q����H����,l���^�pG�(��p��ѻ�IK������b2�
�o|���.��T�&���=��K4 �=�F%+^`���V���7�����55�qT�f�S��Yۉ��e��L��i0�p�H2�l���J�Y�Y�\�۹0�.�6����x'үD�2����ő0��'�9|}oH���u+�+��.Y-ĠK��|�h�b$.���׆�#������U���ŕ���{k��Yu!-����>@���ݍWj�i�����Y�T��l��0y�l�=��������H
�2�7\ē�����~��M�^_���1��T�����QE��ԡN���i+N���f��T���%wT����6��ß� ."�Aw���cfQ�\�b-ٗ1�؜چw����ڦ6`T�f��D4�L
4t���KC�2�	�!�F+��7�����Y�s���J�y$�j'D�^OQ�'Q�/��x@-�-o�o�H3�w�t q�z�Y���߷�S20��suz͜	`��.R�������?�Q�~U���/q�����o�V�<uj��
���*��ig]o��l9׹�����Ӧ���)�>�e�P� ��q��VtE��濗�sԬ��עk7�pڦ��&���e�7�YJ����o���RcJ��doí��J�Ӷ*a�M$z#��)٢�ݹk�;Q?ut&,�<�X���^���T�t��s�P��y�ЪԐ������$n5|WلƯ��ۃTs��7�!*�����K^��5��Q�V�A�Xg�������E����$�_x����<%tx�?��JE��`lҢ���G�t9���-�����u��p/��e�d�Z�Ьa`Y��X?��P��� %�G��2�̪���mӋ{��<?T���^GK��dS$�t� �3|�S����T��kx���)页X\��Aw-��kԂtc�!�~F���݃���.�D�Jns!V&����(�2���Évi$lzT�:��z��j��}$��@�m&���S7K@�Ln�D'Ga���̭�U��#�JΖt%�����i�YJj3���־�- �;���)$O��G�,1lV��+�Yp�ۏ����JncY�	��=Lջ�)#<z�vR������Nd��}�W��T\�"���dm� �ւ��ЏːJ�"��		8X�E���o���ږ=p�,B76o'���L\�B����F�]:�U@���T�Rj�L�2�ԡ�E��5|ȡa��!�*SA�|h��f�w�*�{r�({�8=3x�r��>5����k.�i��0��ͧoF�!V��q{L��&�p�o�ҋe��[�&��Ӿo`��E���)U�:�CK�l�y�٣��dՒ3�b)�YI��،d���ʑ^V���e�"��X��9�Nn�f߹8����{������Ә�4Y�1�&T�[�d�8^D��P��ɀ�>�����h>p@&&ͅ��Ǯ��� A�f�@�c�����[4q=邶�!L�2�a2�)��n���&o��	o�--b��A��.�*q���X�����2ف�7ѥ�Q��+��#a�wf���>�3��%���KH�E��/p����W�J�|r�7�~��B�An�kj�d��8L�n/����u�A�D�4���MG�
�+��y�4y��5VM�
K�D+z���]|{��fZ�^�*���3ǐCl��c�dvi	7��q3J���^��%�&Q���(�qԞ�٣"kn`M���2f���tO&q�C㧩����/� �[�l�y a��Ĵ�W� �jg�>P>��zB���Q�/��%�h�`��^l^2N	���]��3��n��!k$�*&%�����
~��=�	�5� �QA���ܧ��5��q��HK�Du�AL�s���u�V6O^�yS*��d4�+�'�dF\+,1���¿�Ki�*ʮ�'�h�JCL�N�]�<`b�9+�	�苭r��:��o�6͜Y���`��69�D��ß+.�&S:���6�	����u���Gěl)�_��KG.'i$�0�<B�V|\�׋p�x�3L{�q2,<�٭{ҕMj!=�r��"�9U#�,��^�;�X�1Iw�_�v*�� �[�3�E�n�$��*�k޳ؿ�0��8���?��øE"ӊc�8��GG�X�x�}xJ�G��h�:��>/�Q������n���Ey������3�iQ�(]�7up�f��(����\�8���C���/�i,!wQá^����c����R=�lclMej��5�<�Ѡ��G���������]孎*bļ������Z��k�&9_��*�	����KQn���S{��i}�`��Te�o�ylN�5�L�K��ZƳj�Y��j
P[��b5��%���UGl��>�D�Kk�����
�Z� *�:F�J��/>��%{͆���i���c�{�����6�U��j?qcd#O�w�o���L�_��6�0O,�Tb����j�N��Nr�_+D�X���|�l��S��qCIv���b$��e��.�ҐtB��`l�ȭiR��,P��|^b�')X����lzc�>ϣʯ#2��XD�� �v��7��O�ҟ�+ǂW��k�d�b2p� �y2�r	�I蜢�h�A���ax�'U����-��p(68D��jݶ]���hS+��
��Br��Z
��{M�J��*���9�)Ҿ������6�Z?�ߓ��߇��L
��,��qhI\��~�n��G;\:d�뱚G4Zbg�A�kç2P�ص�@��l+,c�z�UyJ��3���U���oMf��C�B~�`�Q���S���Rd#�l�13A��K�n1�[�Ѷs�y�O����\A�d�|�r���.��i�Oً��+�O������M��g��.L/���jAb��tζq,	����3M��fH���� �Hx1��N!ǡ]O����ᓊ޴����	;�|�3��E8���T��?T������W���P�8a	Վ�X	��M��Yf�O�_87�;�<N��7�[����o����=gg�\^ >�ij|��l>�:�i2����(�T9Ҳ��5��b��l>EiA��u������C��s�:n+��x��2�Pt�eq���iy����g��5Q�}��e�}zbN%)��\��2z���>T,q�ߍ�ۍ{8e��:����R�^� Q,B���hF�^�VG�<s���=~�^m���� ���CU��vJ��gV��<F���7�<����or-�6��e�5�?�L��wѴ�m�����2M�H��v^���*����iR��Qj�"�JMiլ���>w�$���B�����0{����Q0��`XƵ�/!ai#07@=5�����
[���y��L�ǅ	E�=N�����r��ȉ��`3���j��Һ�����am�J��*1�y�����\��V_3Ͻ�5XmL�:�T�:n��u�uB����!�^G����n.����7<^+�S�#p
����_���o��Km��|h�؃�<a��C���nE�3�8GVH~V<l���qמ����|e\PrD�_��gkz���q(>�U���d����!g�m,�+�YF��D`#o�)�$������	 _%\���<��A�/s�<�S*a`Q��[�E Q&����Dd�BR�>vGM�j'���q�;٧�α�>n��.�3l���9KL"{��e�:0@��V Z�d"��:|�>�P�\I�̒����A�R�
��A�,[.�9��4�����5��s��Χ�_�V��
�ňd�z���s^G��2EӿA�B���g��ۼMi�8,���&�0�0�l6C�c�a���~4��@�I,�7�+AY(��嫚o�*d���#���%У؞"��#��gsV����f(�AI�%�
��8���|����z᪛1�9�}N���B�Tx���� ;g�%.�&�ݪ>�l\oz���V��>��v���hD���t����ic�0jҸ��
���յ�i��w)2�=�5��&Gt��V;���9<���N�ܫM'v�eQ�aL�K�^"�R�Q�@')u����yF˨��du��nοK4��HK�g��q��DZWƎ��g�� zU7�J��B�U�;hj46���B�R��ԆC�L�O�	-� �q�fyg�l��Xǖ�P3���g4�"���:�@,�^����tG<1�f�\�Z�c�S��&��V)�� �ԣ�Л�'Xv�0�'T��dE�ν�|/�@����1���ǐII ���Jsc_dӎ��P4TQkT�hI�{'�m=+ĜD��7�
�.� g�u�����gl|-i�k�5����'���]p�8܍z^��D�8i����f�D���Q��F*���)gj�2�b��ؑ�Fl��I�͒z�{ eʾ�8&H��6F-������gP-T�o��٘��VN�;O���qhy%��}�0v��p�4]�^@��� ��[qo
�hEA�O��'ãɾ0N���L�S�V36���)L�^����k�\����G�H�b�Ęr�T�����msy����t_|�����L�����zj=Y��}'F,q�.��-��>�����go������ra���j���x��b� �Pz緤ܔ0�.�T�gױA���M��-��E?aw���y����Fюy�@|l�Q�N����%���wn8��~����� 9E*[�����r0,�|,�O7�&�x� �.�C�� CD�����P��.M���X�����Sl؂vpk�EȁA?���-�s��S4��t}Ý��	8�oLޭ������+��GAq�+(c:��(%�h�.��{Q���FpK��Q�%�Zq�P�S�F��s�/�Dx��Wrc�f��L�i�UYs��� je}fC�������i�YI���H{D�a���|�m\#>� �A%�~-|�6|�8��u�a˴�F3a_��.��%�l�~���p�bQ(4��M~�*v3T+��x��}E8�$�E�袩��8�^/b;�P��*��tK�U�~KPlT�l��	���mʓ�8`(�M+�sl�,�!�4��ɂX/���8�������I8�r��u>s
S�ӹ'���Ǳ���=&���
��~�?��B���P��=�uNXL��_��|uz��.��`K�oQ^}\������M-�!Lԛp����*�Y/(�����"�m��1�N�u3�ͼr��&kL�L�ƻ���gO�ϱkd��(��>�L=7�=����q�Xr�{y!��[�y-��ի.����nh��\IpH	�Kzt��k̼~�
�ʢ��#�Џi�����(���z��q�Yi^�6S{ac�.E��\>����	ҶW���}FE814�:,����>::IM�Rk�t����<u������@l�V���k�����&�*{J��UD�[��`2B`��V=A��`5��U{&�/�Ǹ��K"$���B�hfQ|O��y}{�נyBÁğ��1�t2������͌��G<��8�6�O���Êw�qW���R�r=���,��j�p��/��D�?0�'rv���+L���[+P���nAH|:6����A����J&夻m��\��Ir���l���K��*Pw!=��'b��J9r��i��Å}��Hx{9��ïGg�L�=r)bS�fd�C�����&��Jpwu*���h��WG])�?��6݉��-����3I�aTR$Hm4r����t��4=ԠQL�qޫ��Bn.J��ދ���>��k����E�����:�?/	�A�s�#J�5����5�}��Y�կ3�W�|K>8��)H~�Z�u/H�B��g¢R;}l��5}���܄c����>:��ɭb2Dw�䫖�$ʻ�X���������H��Yڴ��+'����r�=��.'���-]�H<
�`����!��l�)v�Z��k��$ToփDQ�S�Q���j�t8_<�t���#X�&���OYp^f�J������6���1{�rm�>�iΗ���3��u	2�?9�>�\�h
=���q��b�Q�l^�d���Ś���o����k�ќ0�`�7<{�V�H=,�PL�Hȃ��F#1�éX �xK&bH��JN�������8JQ�
ǭj�)��lU�s���do��M��]�]pZ��6'�K�:9K~�}ûn��� AE���Z�Q������B�5S�q.
IU��Ү
�E�E����OC��(��X'��&��.=�ǃo��/�d��?h~|�\/����씶��A���P�yu���&�3��
�\����B� ��S�O�4�E�lxp�Q
�� �1�ܟj���a/a�%{�^����!���Ȁ?*��������~�0O��8�}���քw�����1tHlKlKY��BZFR�ɹ�ߑR?�$Fq{� � i������/l�h�k�f����W+��9vn�i��d��h�主��E�ԳG�y1|���V��T����?��|.�.T�䃷ow�\��7X?N�G7�W�@�\�3����vW�E�wӹ#K7��K��38�?��02 a\&�����'B�>���zS��F8k��\vS��{l*U�\h�[q�<��VN5:��In���������뤰%@��3����~]�/&��|�gg�� ���r<�����g]����7Ao}�$�$˥�iEQ��ȝ�0q1O�An�`_u�Z@Γb��ie̸E/�И�F��l�&H��i�؍X_82�˂�J�`T97���'���aY�Gb�~��g�N�o��f�'��hoԬ8h��y�f8ԼF�����"@x 8�4�_�Z���:0w�-H�>L0b������rCwLf���	��~k�5 ��^�RlN�',�����6��W�v�]:vl���4F�Λ�xI�QA9R6�:s�ԣ�VYΚ������ׯ�by�[^�	X�Z�M"_(��}%�!���m-ڟ����8�y�P�/��]8���6�mHVHD3N�X�E��n��tK�7�F.����<Pz9�`&_��`�k��f���ۦй��	�F���M��T9P�;�]�Mx1�l�}�{�ջ1�
��SI�ŜAp��W_T�"�}�r�6�y���A�Z�U��m���ǃ��H.vH�[���`+��:��#�Åׂ~��%�RPԣ������-t���sϟ�p�X�:8j��A]'"~����(����C�.��Z����s��
g�םoE���Jq�Y�����'W��	��ŉVç���� �xCif��+���������*��*w�8��l8hP̃��.F�y���y7C�[=3e��*�>��ݽ�u��|�d����%Q�MKj���!�ca����o�:A��BK^ȭIV�.������Ԓ[7}�\�@���%��+Q����6}S8�zskDOu����f���JR ��& Tm��>+�x�3��Z�� v��z�|}�Y�8��\#	Ҹ�\jCDE��chl܋�U�m�+���ő���|��Jb�@�F=��R�2H�b���3&�ZӸ���DW��ъ�O���k�W�S�[�Se.x�ؤ�J��
JE����N���ơg�43_�mݨ��y�`�.m�Nщ���[�uO��O,�;�X#����24q��13'mu�䌊���V����5/��a�~kS7�u��m*o$|����ɗ�I�Kj����OK'��t�җ]芫,Tp��'���(+�(��/����4H�z�S��Z�}l6�ſsm���J��^+J�|�Y\+��+�c{z@��ڂW���
�M�L���\���
�UM	R�ޔ�d�ֱMT|&<h�XĒ0^a�/��])�^�����(ߐK�cP�Zjfқ��%�;$��'�6�Wh�I,&&2���'���Sȁ�7�X�R���|���:�O��+�G��e!�-I���X���\&���7�'H\��L[F�6���1I$�f�.T.�Oۣ�YN1��������ZBc�/3���_c��3;�+C�#�'��p����o��~������`���G���o��-�Ոl&#�nhŹ����-f��w����#��Y,7�k������0�"���Q�l	�C1A'f��m�7fX#|�H�^|� 4:�
�")ƫ�;�=�����z�U�������\�4 �v�K؁�8���JtI�p�C�|������T8'=SP1B�n>ѮHa���v� 2}��UT��@��Y�;�>*����Q������s�	!	����z� Z�'5�,��	����������������s~R�c�Ͽ�lW4�WԹ�^�g@�;�&F��I���������>�.�������T��K��93�b[�;lR&V]*)���\�c��d��.���"b�ST�(5�ĢJ�|b_�m�x�x��.�d{;1#�C[�����z���T��u���^4�'�pl��<�����k[>2��頉E���]h�ĘÅ,^�X�M��L���������k�c�gk���uMLm`�2ďZ��e宥lץP��=Yi�z���D�Gt
[�Eu(�޶�qW�:S4���\<��`��H���}6ez�����@]��S��8/ *�+�^Ǥ�����?*���s!7]�ܥn��#`�G%{y�+���.j���F���=�Ӝ�O���,�CU 
�I���/m��W�c�I�j�c�A�C�}6�u�n� _;��;���)���>���^��e�[��a����7�AC58�'nh��B+~]^p���윿�֘�f��6r�Xh5�i�f�����MK��B�<u��s�n$�DNd�qR[]���7��}`'����BA;\�IR����V��Z�C�l���Wd�(��/�Ġw{3�=����[3SW6S2�f�p{C��Z�lt�$�󨙽�ճi����<�:����.]���y����ȥ��7�7��m�B�ü������@\F�'�Wݐ�i�"��u�R�ȑ8��|����������g�_l�����G:��fX��߾S��+U'\(�a4��EXR�&�m��<���K���l3�^�Ģsv�������n"�?��>���	d:�O�r�6�����e��1�Z��z�T�[o�*�Ɯ�PB�{���'����v���aC%*}Te��GK;�S�R�+�NR	{�Xd�޻�