��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b����K=&no��|�36�a��o޳�+��T�����p>�����(`W��!�	�������s��?��春;�pmb��t/n��Ј>ֽ�b7���a'��-�B��tl�}%�����ݟ�o(��[�:��<��ۭ
��oP���@�6ZH:�,�g�a�w
��C?�[���E�݆�h��J׸A�jZ�v��z�&Z��ҿ6�0��A0Kj�.�;Y���.}�~~+�7[GQ�C���f��^��������!��eCy>�u�K#��f��ٔ����y��r_���f���� ��ԉ��V�����J%��،p���0!Oт��J��$��vKW�� ��3���,�;<�C�2�$ܤ}����z��#�7�R��J�H�](���B<tY�����HV�4�o����dT3m���~��5:����"�2�Ԅ}���2��h�n;�����0ѷՕYeQ�,�f�}���ϴ���m%��`z�2�wٽyZ]7{�
�}r�Z��A���S?ox!L��7e���}r\�P�4�que�(�w.͓�bm�?}�<�y���z|Ҏ���$}��a������uf��5�#����|{�Ϗ�2g�k^�����w�ex��L��Ek�)�)�G��O˒��F��qV�m/�l=���[�8j��Z�L]1���S����6�����~t��Õib�,O<&N�!H2���=�E��l���W��<9S�K}3��N|b���`���4ՆMM���w6��I3ZT7��(ƼX�څ�zfF�!�����όٵ����[b�"�ȳWή�#�ّO|�^FEs�J�%+���r���T�N��Lw��u������M��!�0>H��妻�����?F��z�);�o+�?�pV�ᴓ�$� ?���!��!:Ī��˼)���!`��5��}+�^\>!����w����60�1Ge��j��(pCU��Z��@���?�){�E���z-K����I���iG����w���e�H	U:��ے�ϔ�(I�0���Fa�GqI�fr�CO5%=���Ь�`�(�\�;�/���FO����l�f��Ë7��Q��ϛ3��l@�a E!������1`�=���%G2<��uo�`�F��A �c9�L��%�p۠�LP�!z��`���Dw��P�^��y�POW9wǤg�၍���Dy���,NW?.������R���o|�0����K#�=��3���L-�y\���t7��ߗA!=�B�S{�kpC5� 8�!Y�(�^��n��9O?oD}P�~�{�s�0:�u|�8����������7&3(�f��W�V��K1�#o�S�(�[|��^꒡��m���^:��R6��W�"�]�E�&��[��zW�yr{Lg
�e �\g; P^����Ӄ�K�!���.����CB����������� ͨ�Iw�_F��5��1p�ߠX��4Ѫ,�����*�FU���5�3�r]����'j}i^>���L|�X��C��>��K��Ξ_c_�Q4b�u���n�_�.�dK�u1�F�P\AoD�N�Tdj^��U��Q.ӎ��;�k��E_�-d�w������ab4
��À~�E�OE�Z!r�9<�'�����l�AW�M���K�;)��ѿV)jf���2�����O�$#4k|-,���/����m0�oq��C��"_��P�up뺟?#]���F�vK:�#\F�V�i�q�I�[�Ё�_ۑELtP��J	2��3��fJ1�J��J�h����O'���Ԟ�!��%�����D���o	 �
T�l�l�����W囼�#��]�����H#��m�n$�/if48��#�(���)�z�UN��2z��&��e&�-jS�����V^n�W1��i�S��� v�D�C#QL0/���σ�j�؆i�����U����zXE��r/��������j��`/����r�h!�I���V �Iḯ�@�tI�d?8���	���"�xFG[<;f���b�d[Z"��;�y	�J�&��>��������N�#�Ӵ��oM��wJ&RU���5فk��c��l;�!�Nr�C�PL�!�)o *��טYy����rް~��i�\EH��1֤T!$��`ˤ�����s(v�T$1	r=T<�>G�&�>��D�k����PN 99�}��T�ȇ�����EMoe[�ţ�=I��Y�OZ�l��86��'bT��ᶣP@���
Kv����]S�񼞚3�����d�\Ӳץ���2j� ޼�k�WH�tIF'�p��d~/|�i�v����MO:f�(��z�x��ddZ�?%DRogM*�b7$9�y�'Y�9Y�d�1
����[�3|$*�d/4�)�f+��R�	�ץ�A���>n鰎?�[0\��'�-��O��i#U�_��2RևA���ת��OI��)�X��l��%��s��}���֒���꾪��\a5�oQKgG����ZN�`����؍x�K�زH���8 l�S��j��,�ׂ��%$�{���v<��ޡ@+\"(��Ca�t"��� ���`K��k��3��D��-9�vZ��TI #��>R�B4�@��|_�b7��e"G����N�������t���,S����V��W�2q���D�$^�k����dAd9 ς.�����9'�*�����)՗�y>~Ԃ�v*j����c�$Huӥ�^Y����3�5���dL��_cHS�]�a���F��B�OM�\�589h�¡���|�����*ud�|�r���J@e����?Q�X����X�k|W�������O)\�3�J��t�	��Ķ��y�[�B�S$N0:�E#S��x���919����Q1���FI�n$�����ʥݍ_ޜ#l+����+� r�8�@!^�ZC2����FN~/����<1ë@+��(�#p�������\b����1���ۯ�����\�U�P����`�q�x+Ȋ˿�rbڙ��Yh�nf����X5��a~d�'�:W��u��G�k�ʉ�C8B�9������z2❀z�$.��*��rOu\��7�����7��0��m����V����ζj����(��8�g������?f����#{6r(�kz@�݂@�����a��(&��&�)���3�#���m��u�ym��0����*d�H�x�ˣ�|>��nT��EV�<3�E`Op���q�{�LT�����{P��g5&n�𾝺;Bc�~{Ĭ����|*~���(�����D�v�Ŕx[�f����]���jD�p-`Q]�@Xj�;-��b`���ɋ����` �<J�ə�]�;p^����1/��(X��Ց8,�Li��6��~��<A����/q)�*��!FX�I�#�(|��io�6������R1�7��[���t����b�]����Xz�FQC"����^�2�2D��r�s�0��]4-B&�-R?�	D�j�sҡ\-�C&i&x�H��PTw�&U�el
Z��r�c��h}�`<��n�'��M�"n#6�\W�Pò:&��b���IQ��	ǽ��E
O�T�zɧ[�ʇ��k�_c��r����K��4� R�������;��lii.j4�yߥ�l�� ��yJU*3Ə4dFec�o��s5����Q�[�������+5�U�g�\;��6��&�u�*�
� HM樈��i����7ʙO\;[�X���.��af$et�Ur7��ʇ̩ �2ҵ��.��ƶ\�"C�C횕��x˺����eȤo�����;G��S��C/b� M��:���g�bnC0�x~,2��C��'oV��uA����g��^\�܌�t?V�/&�99�t���E�m�Sz0�m�P;k�z�:{8���}?/���Xv����6��Vĭgb�W�����)�궙���� 㞆߆�V/��;�B�8�YE���P)r��æ��e�{��=��/��z!��������@�;)��+��J<�����Z��/�i`.�ݍSV������{t�M�}�횯��⤑���Z�t7E��3�Q;��W\b??���:L��� ��Iu���a��S�'qwg�]�Yr�T@TD�7#'@�����!v�����&j�"��FR`��3��#=n�үb� �1��PVZ��>��
q�=�Ƞ,��&f��� ��.Q9f��]3��.
�HIY����@�U����d�8�/�@aȹ��Ws���0�i?�/�L�gN\X* ��	��8d���!�o�D�^X/��h�b��Tʈ��F�8�zs���/h�l:*�&Dַ9�p~�4�"V �o�l��~G��;W�>Ҍ|(*��°��%��s�k�Ў�#��q#�E��~�@��i��섎Ж8��_{D�mA�CE�8(!�6�G�ʄ����Q[��҂v\���
�B�%�{\d�Q�i�c�	�DV�\��9Ɠi����������E����^ gk��c��-��&ZV^�b]J�aXȄ����.��aH'�W�p����"w��4��%"�a��!3�����ٱݝ*���<�U���pwAgF�l�H����V ��r:��^$5T�j�Y]b��ՙ��_�H�Q<ٓN� ��õ��la��o{��}�V6t�w\�-=l\��!tV����F�o΀��I{��ƙ���� j,i`Lkp�*��<G�t_�+
+������}D�4�$~�- #Z��Uq&�ֈ{~D��#�O��E����7~ �n��a�l��*F.����_��%�P�v>�<p��nw��c�U^� ����׵q��2��fw�2r���	�8�f����[�=�) 8E� @	��?T�6@��n������Y�J��
��p>���"L��m��>� ��W�Aߡ4�}�)����������ט߱�HnҖ=��5�	��6S�&}D��tH䱠f�
aT0�3�>�����w�za���Z� �}`�{�L��"�c���H+~�M����7��~*9�6���q�<��yG��*t�S�W�U��.�+F!��-�f$���x���Q%�vͷ�ZtuOl�Y�k�9��Ү��Uq�-�j:�$�1.�Dr-���l��� �{+Yf-KH�6�!�`�H�d5� v��|�AF�/@�ޟjo�|v������a�(�S���++�J�6U ����J(n�
�R��d4��[��7w� �m68I�R�mz�dtɏ��/!�r�~�Ic����L�PӾ�I�ed�J�y�Ƃg���Uޥ���r|�E=�ś��)>�ivt43��1T���-�6L��>����)���z(�W��6�B�ī(ʁ���a�&+S`B;��~B��"_���k�����ϥ�,�~��E����a�tLг]8�1-�{mAI)�U	f����J�1KQ~��e$Po�S?ɍ^ؔ�6=ң߄��H{�#���$ªƗ��)�${on�`����6~(�.L��sW�!*�W���O�^O��3�[�_�D��=t�$1�j���<�����n��ʞzz�����*m��[ޒ���Fm������L)G�0X�W�W�ƊP
�{��d)o�W4��[���&
����[��QwF��Mbe�V��Y��mɗӐmij�W��?��k��o��&B�������ஒ#�e��I�����p�JhD�"\��vQ�W[H�*�l��2 \�LncR�6��O�� ���0��_i^Spuc�^�!x8KO���&.��%c�����Yk�q�N��T�]�I���{w��ق�[�1��N���^ю���,��3�򶜡P���|M��Z��M� n ]���r{LƼ�BbЉ+b[>	<D�z��q��c3%�k�;b2��,*}�_�ܧ��"%��-�P!F%Z��)j��S{��L|��@^!3RB�ꋇ!D����)�|��Z�b�v��]��J�4wx{���b���ڮ�߼xlG_��#�1��l��cU~=���ܐ��nó��,s������[lV0آQ�w���!1�u�Z�L.�9m�����Pot�L�˶$UJZ�JE��ǌ�|��f_�b�L��P�s����Ѹ�I�jBtڟ����Y�����`�f<O�/ovU�xҊ�,�ȯ?[]S�[�p�=��`+�犓A�NY���GIl���q��	�(k˩r��˦�?���X�#7����w��פQ��Um�,n��g� ~NT
8�j��H���=tP�H��`I�R�K&i����b`���fޚl	'�f��4�{�IIA9�9(+a��H�Ͱ�u��>F��,"�o�_6��_eh��Wz�#�]�{�Ϫ:�G��U�����.��u��W�}Yϔ�Gn��Жo?���D��T�U̧x�C<��np�jgQ(��"��dǪj��nMk���$�*�R��X��lJIc�ζ!;�`V�)>�˜��I ��|?G��ǘ/Z���)�{����Њy(��?�3I�ŕ��)UpJEt�������N
�#rf��:�|��ԅ(��y�őP�{�\�(�ď�D91Y1RKMC��u]���t�LVyF�]�}]��K�Pꆲ��&�+�P���ĳ�e��V�%��F�n�5��h<	�;�m#E���K�h��ŉ��%�d�/�1����
J�T>�kj>���"�>h{
&dڸN]�p��i�04��YQT-��$��r�\E��F��#�.\����q�$74C��@����s�1���d�a � ����.#K+�<����$+S%����-Gu�f�;�(�NJ^�F}`LjtZ�ש�G��s�GR�+���sLM�)O4���:�Y1����eƷZ.ՍڌڬMk�ºB����������!��_�B@+֪�Q�_�� H+���P>8R�u{�;�>ټ493Q��0>27剺}�$Է[�'ACM&�dX@4@" ��^��ƺ*�����+B����RL�����"��f' ��&����)� #F�Al��F�}%yē9u9�J�9�|#�1`�ۗ�]��S�fv為A�hWWpʣS��������v�����i���п�p0F�$�R"E��P'RBM�r�uS��1�ￔձ��/z���>��98��b�IL| ����"���"U�A�[O�zu�zE�M�y*���g��阶�f�w��dAv[O[C���ܝA��'ry���ǒ�&������N��,w+d�x��[dR���ZX����?lI-��,��wAy�d����FF�}�1�y	��NT�����}.��pu���杷I�,�\Ԑ��cA;��m����P�� �|�~�=hE�&��.
	�9�:��'R��C�N�rLY�Dm�q��D�5�S�.:��|�c�y�A U4^[pU��2C�*�O�����@P0�#{��ݘT��"�M��05�@���4ބ�t�(����}v�{���g�y�V�R6��N�=�7�"}�GڹB�- ���n�{6Ur�Ǐm��&�SR>�z���i�LI>�U�hY�`��\U@J�iEL>`�
Y$&��_��#�8�����K�l�lWu�7�q�l��QqB	ĢyCmI<}���ݔ*�f�l�����MSmS@���k}�I����*��&4�	a#%^螔�q=SѨΈx���n���B�Ȟ���4��8!�%��L�c�Z��4p��O
<�;q4��~�h������@*��g��/8���h��/c�,�Y�6��q����{�����{�J�`�k���'����љ�	B��C�'��-pS���$���0t� ���8��o���j4�u�/Cb嬷���9�c҆8��|w�K���-���%%���z�b	���)e�n��H�M����V���M�VW�d��#pF�r$�_��X��OӢJCVa]=1�iM��UR���E�K�2+����Pz7A����GDwh|�`��(��}��w g��
g��l�+/�:�����a[$]%�P*�Lcty%�����1g�&�n��S@T�,ۂ`�����wd����2�f�u��t�@�nҊBX�Y���O�����C�Rjm�'���1-�v
%B�'�mÖ��HG�ۧy�k��グ����ೌ69b�n��}˓��р��(�*� ;�ğ�Z��<K!�3�c��0�-zK�N:W�>wb�:�b�R��}ZEH��$|�2~�y~Zגuڀ���������W>��r��r�.;R,n��h����1�tIC�&�K�����:�A�b�\P�kw�iM&��ƭ�¨�vc�0��a@RAϭ�P�����P�_���A��EL�-a���?зM�\�T��R.�.���"-������qlN�Ɉ����w�M�T�GV�M��c;J=k����Z���}*�؟�[R^/�X��?��w��z��r��^���{�S���:O�p̀9�3��[���JG����`"`�BÎ�[d&B�M]E��>d�������&��#/]�;�U5�"'a#�g�8W �9����tϦx�\��ʓ�@����Nէ�a+�*���PUDɺuK��]X���e���|��yPNk���m��H�ut�'����un�v'�1����?�eb�z`pc둘�U-����+������z�rSy�Q)�������H; �6M� 1qk�'�N*���RY�[�ֺ	��Sѻ�S�ʰ ��(�Z
Yh]�W|�����n���9����M��B$$E�.V��c�;f�'�8�B�.Ơ��#���GT���续%��*ͣ�W�N��q���E�S#.СrK}�G�}P��AP9&����&F���〸|;f�E��B�z|H�2��O
�i��Ƚt*L�0�B��\ɥs�;����}q�3��1�,�����)�qA�u��OFi��~@ɐ�	H�zy �@~��b�.�n��;Ǧ���}�:�Y�cl�JO�q�!s5^�m��
F�n�������׶zI�|l�a�/{d����?��f��O~l�b	�6�T��.�Z	�E�c@�W�&l����i�cV˪�o�>�+/8��z��%�k#20��t?=�)��W�no`����π�XB��}���n��d��H��w� �7�<o���(7�� Vʹ�W
))S���2�yfQ�4�R���R΢����9�֯�{�&$�͘k�R���S3�j�.�E�zֿoC[����/<������ˑ���\/�Cz7� $�@h�Ѵ�������s�&�It��J�����Ǆ#�}q��C��R�,�ӘW�s���gt��M_e˚O@A�̋j-ݿ ��C��39�{Z�uP~N�g}� ~"��*�x�@u���ιW��w�*b��|l��"�qg��|Ui�p�նw��zG�7�>|�����1i�<l�"�A�`�? ;�q�L�(Ѵ��a�m�u����s�K��8{�MD� �VĘɮ�}��}8u�[�Dl�e ����3��hI��u�׌��LO��5�����d���^id䔁"����Zē�8!j5��rR9��,�`�睅�qE-Lfʠ�m��Ĕve�kE,IU���"��*��(����=�6X(R��XNM׼]C�b��x��L��ܧ^����wM���g�X5���}C[#�I�%��5!P!<s�����7�PTF�2U�o.�"��Wb=���/���*�Eģ�$R&:��L#��ۿpʫG;<Q�h�2��n+yT�?�:!��W/2]B�����HE�q���{6Y����|�CK��v�R���s�!����
/�a������q�P�#P}���d���1������]^����������l��s��������p�u�N�]$�'N!�t�m	5(Oy�}uR�ㄌ[�����}u�9��S���y(Q�S�X�#1�Ҏ7��W4��16���E���AXو�l�1�A�Zh(��3ڷ��!�2�R
�PaH�I��R��	]_r�W�,�@��vu�����L�a���}Y��ԎC�e4�c�ro��/*kh�(8�{~!������4x� �牻��*�_�Z)!�g$0���Q��zϽ�ɓ��j�����8����g��	!�Xj�C��i Q��h�^������Xɢ�>a��ܑMl+Ld����>8�;ly2|�h���=�*�P� ����W])��y��<`�\-/�Т�S�Lu�u��u��u��%m�h
m�{?9��c:M�"���m[�Z8OY�c������q�/&}MV*3q��;X7�lJ�m���P`��H�<�C�d@%�U=�N�B-=���u�=��ިo�e>8<���=�oe�-Շ�wY0��D�0�`]��B4��E�'c@ѯ��*���LIC���F�sW�NK<ۑ�����6�dA��l)ɠq�&�?pv��=�(��]3�����|e����	�_�:M-T��zsF|�Tz�)&�"ۢˬ���f�
�ú�x1�|#��i>���M+�
.^'������� ��v�TveD�%1 ��^O�6�p�oib�*�Ys)�:I�*�z���X�f�z���EҾ�.���מ�����Q����M�]1���/ɰ��ؚY$g�}���`j��im�k�/z,����g���C��R�WgAj��o��ԋ�	]�1�R�X���+V�|�|릊A&�=%]n͘����=��T���"7��ת2�du����\��$.�u���/Ɨ-��u�� "ձL�	�y�1�ͿͼY+��	���]g�\�܏�^T����2��P*dZ�b�j�j�U"Q�ܖ���y �ڰf�"ӯЁW�1Z@yc���W`�C1��H�O�d��A�:U����z�]���[��k��F8��/�����E}��k#-tn�+$�����k��mÂ[T��)m,3]�u�Jt��*��2WGPGM���m>'0<5#��(��/:�̛+3M��&�ك�P���>�Q��W?C�[DŶڻyI��6z�XT�><�]�������01w���INS����o�teF���Ch>)��J;LS��Z�j��o/�4��'a��*;�h��C�K��3G��r�p6�L�vEg�~�Yl��ԒT�j6*��%��y��jv�kL�+[;�AE�h�F;��nݕ��ܽ�����Ssco�j�!J$�m�R��jng��_i�+�9Ý�G�|�{PH��>�_���{�\Tl��`�t����� ��izc��x�)�P��q	� �3Ԋ:��3E#ys�T�Y�<�^A���r��O�~�z\b��3x�ōJ�%rB�K���d�� �C�>=Ko�W�C�z�������e5pnS�7���@I��U��oO�	��h�B��tl $�i�� s��#Y�hL�N��w�dW���Zܕ�rZ��	?�`�EA��xN�J�|�u
j	�Ȯ}��r?G�����o4��N6o6��a�L	08π^��]�?3oML/<�hN[8 L���2*�k�9�j���c��,��4Z\,6a�ze�?�A�52d6���n!�(�}���1��~´�TA_�lY>���.�����}5�$��"s�1\@�:Z�U��N՟ިn9HY����Rɶ-f��x\���EG4G�V�R�(qDΒ
n��|��NS�����a����
G�X�(��|��5��]&�溥��)�����ʽ�L$�PbwC>���<���@�1�oGJ�O#"��l�	(�U=�Q�i�!�=�q3S��Y���g}�:�s-��[������RC�S����	�8��>k�Q��!1e���SƸfFe%��f'7��r mڼ���j��X4k�:���>C��(��pԶs*�G�o����U&��0½ �*t��X� j����\�ȴO�V�'.�eq�����6X#@�v��L��\�����9'K���uBu��q��&F����w�pЍ+���@k��p^::Ty�r���sl�.�8��s?�w\y�n~V�R�$�9�;a��$��z�����?T��l�� y�0ZCY�&�2Xn���髐4����i�eB��IjŽ)/0 ~�����:�2r���D���-Q���[9&/���` ?�B�K���ZN��A�Ze�f=R����5zޙ$�Q�5o���-�5'�*���.����1p�Z�;^v�}vj4پ]����[�\�^����1^{Ej9h�$�sl�X!��u?�&�J�B�u߹o����z��ئ�j-������V=����_��f��%r�g�r�1�=U640_�9����;��֠p���liz�	��	�xG� 8������,��z' ��
�TU3��1BHn�M��38����L�E��= ����)�ޱZ��K�\h�H����,Yn:����ܫo�3�Op���BX~���[�D�M��2���3!NX�m�O!w�pGw������ہ��p$O�㒄vZF@t��53kE�xk�I��,VL_.��������k�_Ak�i=��V�*���UN�ZU|گ-z*;��L�$>�R�a[�M�[�V�QTp��s\a���P	�	�Bם�m��*"�xQ����^$͏������_,���L�@����?���9�T�h4À2��m�)�p�v���u3?��G
�)ޣ�%8�D�3�e髞U��q�_�a��ugN�wj���-;y�}�����r>��r��_�~Ш���ު����gf������}ᧄi�^��D|�pNS@���YRL[կ^Q�|�Y@�I4I��:���N�0�@N��$�g�`Q+����R�)Li^�)�P��@��/F�1�j��I�:��Em�8~�
Naբ�FN�{/�v���[R?@Pj�[`��.Pz�ӳ\1�����(L7�xp*rDatOp.K��b~�t�?p�~�w��0����Q&j�͋	�u�5eC��Q�Ƨ��\:�:N%Lk�ľ�2����d5�?{�U���oJ���a�y��� h�>���$��@c���"�J*p�:�u�@��Rsw��!����E�O�6M����-��X^S����o�r$�ɘD:��2tC�/E:"t�)�A��s��S�Zy,��^���i��
K{f�h+�	���(%�?g�J�^X�9�b�g&=��������s��	�f�Y��C �$ͣ}3�(C.eC�	#����^��a�3"�:���H���.��.�����K�~�$��l/Ŷ`�.��8Puey��䱗��ܮ�-Z�@,�~<�r=�jB��4�e@�[4_U��h���/޷���4o�
qS�P���Mw�Jz�7c��o6�٥�! z��+5?�hL& =��*��PB���]?���1L�����������d���s