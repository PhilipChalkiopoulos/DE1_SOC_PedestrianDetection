��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���jl�7�x�֫����_��aoY��?#��#�r�m�"R^F�(hb=��pt$��e[5�v� ��n{L�x����o�x�+@wM�ca冐堏����D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�NX�0A�J5�02ye3��<�a ��j>��B�q3������h@�J��f��)�d��f���-�!D���xv/�b��+���~�q}S���x�g'n�F9g\��3�O}�L<�@�G#���$$K��w�P�6��2I�ޕd")�W��Ғ|�!0Bmx����DC��%95��X +��,J�[�t�/5͜���?*@'���m_)�M���O��1�Wm�/������c�+��0�,�d8�ŭ�ׁ����~(��m',5�=,fRh@4kG��.�N��A�M�c)p�(�B���&�{��Wi��@m،F�|�����*WqBl���=��@_���[nH캺����]p&����19Px:�5�^)Qlo��%� E��7}�4�� �B�SӅ7��`$�����|����w¬�M\~G.���ړٞx�_0���PLY#<�̦����p��} ����ܕ׾�lM+y��Vb,F��ڃ��}��2���J�	lr^���Yaߦ"Ţ�`sFD�Sv]Vܾ&�����_2g���-�A�tuJɣ��L�R���n_ֱ�	-0B๏��>�ɋYq="�+��qb!�X.�O M6���@�9M!�2���[��!Ex1���f�m&�2[��F���D�>���L.���«����n�oS2��Ǎ�e��[��p՟���W8��W��C��9z2�������l�cE�a�A~f�A�\����eU��3��7�QI�J����|�~�Pv�fPq���M��̂EI�p>���޳�4;�������?�c�GC��"�G$�]�%ڸ�"����ԞOu6s��n̨1����i��4[�9�2wOw�U�@��l�� ��c"��ي�y��U�P���Y�:��4!.�r��������B��A7�y��?>�$��0��s���;R�K��LS��GcG69a���Q�JF��nD�%i����qwǔ�kJs���������?֩��_��Vp��6[1�v��ԭ�K����n�@$ ��h�Bݘ[�G ��
�a������ԅG�ܿ�����HǶ}��ȝGS�j�&�� )6yej����*�=�����������WW)�<р�e�1��6
�rfJ����4�eU�P�*��0LZx�][u���h��͕�j�4ܪfZOE�o~�$3g�S��I^n�ݬ�f��N��K+.)��C!��5B\x7.���;��f�2���Pp���x|zڀN՞`�풂�J��H���!����X'g���[5ʾ{�U{�����Q�)��k�
��ɢ�2b)��F{S"ѭR�&U!�*8��7�J	����o*:��5�]�2�vL&Fx%թ���Z��l?�o+X�u��Du���4���Z�o�V���$�Z�"��67�1\�(	+l��9uC�B��UepÙ�Ya>��">�nZ�m㧾�إ�₨ڀ8:x�Ȩ���%8Tz�-����8����+T����LYW�ț~�q`[v����ܤ2��E��c]��R}䜅=��挦�͈����~%��l:
���e�S�t��mR~J�Ĩ�e�9�P������[�Fv��^\|L|�钦[p&r��
\��E~Ls��}�\�}a�S\/�f������ 	�oV�O�m]�(��Or!j=�ȝ�8���9Y_ܳxq	��b� MEq�t���~H��������	8���Ŏ��2����j�FOO�(Sm��Z3���p�f�{�؎˪�^hʬ&o�D��{	�����
�t��Bfo�YK��vv�mWm��S*�ݶ��2&�wG��[���]F�9��!�}�Z��Fb��QAr��Yy��y�ke�O� �k��J:�=/%v�F��}�A_��?�R�R���!�y�vTKH5�f�k����|��p�oN�����@�B�/Rz�s	��)��#�W��x5�� Y�s��U->�q�G��'}���k,_Gm�,5�D!C����GZ �$�5��|��Cϗk���;��N@�lB��W�Ъ��-��4�L�����]nB�9
 cD�X��������ؓ��oW|��ں�d�Em[(jCO�; �W��o�
w���G���f���!�m��蚣o��m�����ƣ��"��=�"��^� �.%�iO��?������;�r��S��3�P��\���g;�
�s�,R��;8A��	�Ō�s|�u¾'��z�aǱ��� �=4k�������	�Z������b,9�L����b�f�+���)�p�����t�sk�L�7����j�L����޺l���=����)Ir}\,���W���X�#��vD���}l���p��$B�_"�υ��=�a�1m$L,%j|��M"�g�v��'u򈞹=�y�4}ئ�$g����SF��q& �Wp���v�Ÿ�l������:���Z��o��BJE��U97eC�:�pH7b���q��rTZt��Ä�ݰ��H��FWŝ�w�a6q��WA�I	���7�T���y*i��NG����|<ks�l��D�,́��I !/���l�'v��^���K+�
�|`�V���0<�R��^fu��L������ܣ�d�`NE���H�!������?�G �$�"�!f����%�ܗB,�v��e�:�N�~�v�p��������ľ�"�^�XEl��ݗӋC��jŇ(R�i��gØ�WF��I"�枩�=h��~%l�2�1t��Ǽ�}u�ƙ&\��9���R��4��!�,�¹!�;5��ӊ�#6��b96^Z{�0J���x��^M�mf��G�� ����j-L�������Y�:�(<;��QC�0����0p��C��� H�A�'�S6!jo����1���o�r^��GhH�[K	>JS�ma��`��0/�a������kG't�{Z���`�)Ӻ���x?�&k6�%:h������eϱ�7�Zd�`��l�����i��|�x5~o�2�Wjq�u6��;�O�B
��������L�>�N�}��SI�@y��3�q��V?��>���)-E����aMvC<��&�2�2C1���fS���K����9|g��f0(:��v������_r����_����y�*�9��PCߎ��zI�\1������{�e���z�vhA{�p	ټ>w����kK�*J&��"�	���$b����a��4��� ��n�_�tw��K�M������M��X�>�AY�1Rw3>F�y:�WP��<Y��𽵬�@�ň�������g����Ê�9�o����v�\��~���/�`6M��,X7��lm��� �my�ґH�Z3c��*�m�p�$�#*�&W<L,d_r��N|�������L���y:u���f����:�I��4��5�2�G�Ӳ�qR<"��"K���ܗd�p��H�4�H	0#��Z�!g�(-J.��dС��*o�;��_0����2I9�Z�=�]}�.���CV˥<A~��Ǔ���;����Ⲍsu��PN��èe)���HPKB����Ȱ�ay�8��>� ��m���J@�ST�<G���Pe�r��U�] ���Uy��38s�&��l'g}P'4zI��Ma�ʮ�'^�&��k6��b�+}��|�D�fU�Uq��Wx֮�lݢcUe�o�St����6k0S�]s��q��@w*ǱN���� �ErP�`��jgg}���;�j��"����mX%�(�7��-�ira�o����~�쒍�H��a����zL��eu�c�W�j| <���.�ڦ)�k^�crMI�D�\�bgZ��<�������Z�<<ϥ��d�V9C�����b��W�s	�yb�\��\1<���ˉ�E�*j�yMٖL<�>��]�hh���O����Ǣ��=�c�r?x\��Z��Aв�.�O���⻾[���}(L�����-3���IF�d�	U�gx~h����[y��q�;.�W�ò�ɵ�6�-&����k�ኆ)�P��
P�.�ʍ6��P[mvR�.�����l��q�.����V�uGբ��j���Q��yr/���DA�g���ڄ�W1�h��3�4 [�M=�������.�,����}�/�y���gl�7qcYf�Q���	c9f�5��Ȫ	��>]�X�*�!r���X9�0�xr VQ��Y(�^~�8`�7��E�f��Ō��6'zI��Y�\c܁ {������+RY�N���B��>��k�0��1�ď������u�3����&�3=^h)C�h��5�'�d]QY:S�S��"��9s�X֕�N���&��>������zz�|q��-q@��:b�	G��$m�Y�6����b#��_��X��%4��l���c����o\������j�>��5˃��<��w�ƕs�Lb?��m57}��1����=73�*wܐ�)��봯$��Q		�Ũ���Q�+�R�t���q%�^̀��K&�b�)��z�M_g��]V5�%w��ʦ+g�[W@�]s���%�{̠��������4�l܄��[`�S��]�Z�:������Y�$,��ք�����ZE��M2R�ώ�����,�A|�m���S�ܰ�a�^�d侇����B�1 ��6ug�F��_<M���,&K������0"+���-l��Œ�2q����25f��-���:��[Z�P� �bۭ����ZX:��o����VcVZ"0�VH	;glf���E��yxCu<qJ�:��^AOQ[�bh9�h@CX�8䕎·+�����5�Lc���X��Bw���LX$�*��(/%�,��	Is�I�!=AAv����bb�8_Jlz_��Dl��;��L]-Sy�[��`�H��j�ջd���͌����}�Hl^R�/��+���m�s�&�R���=yjw�]4&"����G �R��G��׿ ����ZmZ�����8K�my|��Fs�'7ݟP$`����\�mH ��B�a�1��*{�T�k�����7�En��������+Pam��{� ��U�}e�p�!�����Z,4�j��
��ԕv�v��'��;�ʆ�@~�#n��x�c�Y�E��=$qS>)3���n�?=&/�>� T<~2�2(E���Ϣ6��8�&?�vQo{y��$�h�b=��P��EH-��[J��%���gd��y.�"�n�4%r~�X��]�Kb����ۤ�Ⱦd�'b`�T��4́ƃ_�������AB>�7�$Ɗ�,Ya>��k�N��)b=�y��� 7��:�9�B�al%B��dI1xh���WW�3a���-1;ZaX$��@�+0�B�ݾ�����$ލ�⦬���O�z�#��*��/�(���v�C��*j){5�a[�]n��'��xVs���%;�zZi�7�<(;^�!�_�����'=�!VHO�'l�
@H�u� ��ٿj�w����]j����X�32�-Xa`�Id�X�UY�&���&�Sli)��R�`\{���gV}XP:��?�6��%O���aʷFVNj��f���YN8��D�.Ȱ����=�X'=ǜtb����Ʌn��KU񡡉�LN��GND��ڐn�>A�I�m�W�o_�����ޠ��[8F�Ǫ6��@C�b�A��ݙ�_��i?Q�����:X�c�1
�MDl�[0�t��ȉ1#t�;ޔ�a�|���y�/t`���C��D��Fr��;��z�����O���[(J��˥ T�����I�c�����I�Kg��6��k;ߨ~WyE#���D#<�%��:pZq�/� 镏�_��SEJ� ����[H�/ڳ���m�fm��u�㦉�I����Oѭ��Z`#0���䚂֖2�qo���|r��╢��ƚ��\�8w�ԉZ/wT��5��ki�q���3��f1xG�>�!)��f�z&�#���g_o�N�b�v�DR����m�����]º����Qi����L�ʥ�_��ڀˋ����3W��������0�f=�&蝮�(�B��ppq24f"T�dl��'/G�t���+�`(#�*>c�y�%#�T;����S$��6N�7/	��գ%�F��!�4�ԇM���l�b4�Eu=�G&��օy=[U���'�r�g�W��]
���Y�����nt

%*�u�WCċ},f��.��}ߓK�if��ݿ��q��t���lӴ�62�6({I�����D(}�)���{��7�M�}R2Fr,�����C8ַ^�=�I��dWĿ~S���^߃��LfaMY?_�G�C�n�_T ���
�i��R�Y%��o�;x��(@��f��=U��l?+�f=9�����i�d�b�_�l��8�Lȹ��5�{���!��x=�;܆*���SH��)]�g|��*՚��b�[�Gͪ����c�"˳��q/im%�OX�o��\8��7 ��ĂR���W�mǋ��>N��?�gÖ��c^�k�|D�=�/�6"�v\/1�����`�d�����D�������.�v�^��î/"'J��үb�S�.��:'T�k,����I�ŌoK[\�X����/��1N���E0����z�6*��'�y�wqWݾ��J���B�IY EFµ؀���v�cz6ک��S�U�N�h'��5�Hx&&bz~���I�5�8���e��3���B�n14eJ�lrLs��n���ۯ��3;N�i�ㅽ��Z����l��U�7>n��s��d�(P����Q���H�%�U���2�:ɕ�O��T�#�B��K��e���aDv4�����dw���Ncp�uhT @D�X!ci�E#2r��0Q�'�s�  �_97�j����$,7v39��sz^�p��7~dA͚���r�K�P��\����e�b�Y��� ��(P��߈=�@p������2���~����{�v�̐�O������}.#���N��O?Z���~$�l��.;;E�U�B�ӥF3.$�XŅ���5"�=2cj&*���~�c��j�5�[o��ye�ź!L����|8~q�P�;]�L��ټ��硭���6�\q�ɓD&���F�Me��t�{|��F5xV�A�Y��^yס �paz����H�s�z���*ts��k�''vۨ�c��'����1�X�Ax ��
j�o{n����R��u��O!^j��53FQ�s�����uh.��F�+��Ve�aA�FQ�m3�A�dU��|t��|Ç�� ��|���)��ĭ���g�y��>2��Beޙ��*�2`z���q#R+�@�3M!���R����=�L�v�(4�v
w�s����ZR3���+�1q�'![�cPa6���8[�Gm�����[ۋ��F����C�G�V&M\	���k�_�x��G|���%=	7�E$�Ae��|qׯ��c+>�_9�r*�	V�v^�}�R�sy�c�_�0ι;� 6�Dlt������b�WQ�wڦ��i��ӏ��q��Uմ���]�I}������<�u�v$�l�<<��h:��^~��g�G ��,���h��Y�R>����K�����+ȟY���+[�Z1�0.� ��a��rL�XfJ:?�DFH�Tè�U
kpY���☉��r�NTs�T��,��WBU�R��s�FI*��:��G�Ζ��D�ٶW�U�����4�/���^�Χ
��6x���Wp���:aÕ��@�Y#�|���+0.m��t�>���5�
��@���L�(d���(x	��Z�V��N?���wI�瑣��s��\)}�`����&�J۷-��T����g��j����g���.N&Y�T�7-R��d�m��25�n&����re�aF��D�w;�k�~������̐��6[Ea6�O�D/0̻��(�F3���=,hu���a�	�Aګ�g2�Fb^
G
��Le#5V�X���B��23��wD���2��Z/���TC�l�F9�������GV�SAȠ/�.X�?��2�2�f�����$;�\��¶Z�5�3H�:ĩ���3'��| ��\U����c��*�zh��	�R~��o�w��g�x�\q�1����ͤ�
&Y��[�@�3w����߰y|O
��D;��/�[+ϙx-��h�!��kG�B@!1��ߦ I�����sM��,R����>�O��f��H�4O�T.��� N
�d� .#�p�`�q���<h�����L_Df6m�{�����J��`���_p�I�Պ� Pԫ	�)8.���r<j�军�膱N�1�o�ы���¾u��Y۱}�eݨ[9��↹Hb}eϒód����*��zt���ҝKߘ�����5+�l���J{4eO���cǃ�0%!�L��0��tq��j�:|h�]v��:���d�/�>�ع+�l���V�bp��2�U��%(o<���]mc��c� �[��J�����%:#�U�ď]��VM�A�X`5,@��O�PJN��;*B�s�j�0nS�� ��l�k�v��=��_�p1#cT̸];�Өjd�4ٳ#�4�C�h*0aL��"A�,\�����&�dSǋ��H���?5�.�Fƒ*����_��������y*�xq����
K���TؙuY�=�����P|�\�q��^k��kG�6����H<gM2r�`5hye�_�$X��sLe*Q����p�������y��d4Y�����PU�f��m|��Ll�@:��c*+��wp������}_�[UP?Ƴ>��j��|��,v{!�0�ڼ�mgs�����P�z�D8xͦ���D���(}_3
���P"3]��4����=M�1�V
/�8��yX�r���F�4�_R����B�u	��o*X���_�pM?�p@�䵸�h�&�DlAa8�GVbU�+���W�N<�x�+K��:����Dƴ������'��p�>�U�n���p^�D{Nj�H��q
}ͼ�Z���g�Ni�r]�����G㝫�LV�pa�*�ܘ5��:D��K)�; �lᤏr����*�&M���-�����;U�S5��C��xP���F���P]��lw\Y��ж�)dփA�v�ڏ˫�ZI#���˝9I�B�Iu��^�	�Ҡ��x���c����0��d�r�8�:)�f�-9/���K�x�R�-���`��2�s�&�b⑛jkd�sX�S�s�����R���	1t��KA2�fF�֤UK��;q[�u��:�U�y�u�:O�{�%�e��]��SEb�k\�;�y��i�oh�>CV�]9�Y�(e�<�iON�i��~��[�%����y?|�9����L �f�j]�z�������1��!���q1���Һ�r��,��,�f����B����m���Wk+.5�4ZLl�z�Z�t�+,$o}�6�����m�T�@�&�pm�j}l�&ԔRcCN���뢪��d��r���L@�R/(+�����ȉ�ɝG���|D9d-���������@�{�;+QA��S�x4�j��aK�79�2�#[�u��]u��{9m�MU���^[ �{�Oޡ����xG�]���F%�r)7�0�:^������w�)�Z�O"���W��2�h/�K-��%*�k���NC��������<�Ra�Y��b�>�kqF� �d���WR=��*��[��P�H�1%\o�$.�3���P�P��I~��uA�X']J�B��7��A��A��&4��FO��!�{S̨� %5ƞ��W��;#��0��\Q5`�x\e�}k7�'|Eč���(e�'��@U�Pk��JI�Q$c�Q h��T�N7��el�Y�ₜʻ��U�Y��	JB�G�Xg�)���ji��Ѹ��i5a!�[dN�=a[:*��n}�*�W("��!��~P{�D���d�!�2����%*���)�C=��b/.��%B����jO����qpM���sws�8t\_��m���+�VP�wH��]a�ί�H���@D<΀$�ϣ\ i�&c����;������-��N�]]�I(&?u��RM��	���,��p$&���b�م/H�O2M�5�Z?/���%�9��:��I��7r�O6Q�:�`�?���dS636Y�N�j��CuWq�[ز�Na�9`� =���%W[y�{�Wrˠܜ	Lu��7Y�q]Y3�N#ȯ,oI� r�J���IT�c��p]{P�q4��X��Q��},)Fx0�y�x�X��x�r`�U�؍D~L�.��1W�Re k.h��2�M���ܿ<g|�|�F��C��T#�߶�\�+ܰ����L��d\�������x�Z��3�@XЂ����>r}�~�
N����Z���2��{�@���Q��o���Y�A�x.���:"z�刾�'����V�Y:���r�E��27�w{|Eşg!�ƺ~�5>>������O\v����f>��ο��5�W����.p���8�"����lA3�F�N�F#�n:O�$yFc�u��"�:��d?�B=��'�q��I�1:�R\�4����r�2�IPz[�2kzP}����;�Ȗ%j�a"�BXdC2�m?��I��qW9x�*̎�*�rwOk�B����>GZ�ed�@����U����*��n��l�~]$�6�bV�&�l�y!|���M5<ɸUfC����*@�
�l�D�)�\���ݾ��`T�w���w_�����TϾ?F�������ȹ�Wa���*<%j�u�}�}�E��Bt@a|�ĢD5�8 �f���1�����LC�~?�mɊ��3.,���*
!+�����<u�=}��_��b�N� �i�����+���p��3��e����(�H4�?��e��Z褪�VAO��ħeDސ����'3����(��\�at��'Ì�����%mѲ��F-n����Y�����餐͂�̻�݄v�`��wZ�*�/�����
5^�I�c���S֣����3�fo҂=�,|t���������JJn�A��"�&��SU��V��$�k�d�_�C�5,�&��*��<��}�OC\�WW��@�ݺ�I���k������m���-����[��[�>�H��� �� SYδ[�?���8��ǲ��Pm,Uz��y�*a�/_�D��?v>t�Ƴ�������OV��Ţ/�g�O9�j�Z=�[�?G9��z*�A/B�Zl��>z�p\�i,�wY-f��Ŏ"�5�"�k��R76�iP0��o^�P�0��邡.�|��>�&Rw�5�]2� �l�"�#�r��&!�y[��uTW�	̹�oe�\�蜂��`L5�J��p5a��|��~#v�.EN���i'<��Е�ac �*���h��ɦ��i��s;ՅWmb�޶���=�"p���5��J���^O���A��8���o�e�A��ڐ�"�W��4��\�ިN�{��8��T��I�����&��+ ��j��N�^i%z�bGV�D)�/DtT��{s�ٜ#�n|�'Ҕ�А���������<��ϴt����#@�3��-�'3��f�sxg���Nbbs�P�����`z>��T7�(���w�FEs�P�M� ��G�)x���*+37�p�"S��⬼>��=W�,�s"�q����k(ᩋ�f�i{�k��Qڑ��'ms�(��g��:�1�Ǻ����/K�Ц�e�ӗ�'�h��ˊ.�g��F�w᪠�O��=�z�2 �U����f��Μ��d����0�*fo��$t�}w�}}o�C�F�,�+\�B)>�[�����%�Ƒ��&�ayv.8p�i��DP��vK����$9fD�;7V��\�RفJFH��d��R��V�>��9Օ�r�KL�{�k��5�`�~s��"����q�(�Ck�o�O�F��%��3V�
��^�X���x�����􉗢�^מ�� i&�X#,Ar���V,J��F?¡��z��L�: ������@�6S��w����\�^^��R�/�3����z��t��I5>t����X_����wi"QO�lpb�l���D��e|�g��p��i#P���p"]�R�uyR����{7(:�	�����/귐$�3�
�E����g�]��T��d�SL���gFE=��"���.o�c��J�N�*����#gR�,��o%Y'�O�2��f�aO�7N��&H!���:ߊ�+eG��'Y�%A-�׎�B�� �%���ȤL>q%��ԨH]��5�n7w��M��Zk��=hsz��
�,ˤ����/��-��-&�w��%�v�[���y�D4O�`g�v0�ək>�O��r{�1�p�D.��~�a�k��T��b.X(�7N���?u�GҊ�l��3׿�K����@�<��y�yA���4�{�%T��+v�k,��9�"��LeJ[��������0�~"=��Vpp��h�`��U��e�nWvtd�0ڑw�>K3�qn�DQ���"�[��l> ����Tpb����\�\���tZ��!��4���"A�3ym�c��J�N|y�^�����E+M꯾3�i���K��|-1o�B�Wl@�yݬ���ꑯ� SA��m<�A�����D��M*;�>	dA3ض	`9ʭ�f�?e��G��}��gd:��O��R���KKc j�""5y�(�CvAvE^I�1�7�����2$WŲz��T*�����W�L��n ��T�p��j:�X+0i�o�h]�]��[/��˘�D����r�n���m�����Q�3�!�:�4}7D�ς��3v�3q;}#yu�>	z�[F9�y�h{�:�x*�X�Bp���0�[;X�NЌM�ns7��>|���c���E��g���XF��F��2��+ٞ��?�b��H�¸�]K!W�T����Is.��c,|9�(A�n.�;H�p��9�#����m�dsԕ��6�i*��1�� ��"�����:�|�� &�c�٧�'�ߕ��9����e*����l*��{��;�(#�D����ۓw���������N�f�?1���%�h[���\��o¹ ����iR�c�����r���Ǘ�^5dJ�Dʡ�ܧ�n�A��7���Z6�`� M�=�j����zu��1��S��&Քl'��W�jx�L�@^*¥q�1���mm�b��YMu>�,�8BZĲ0P�bZ�g�R������{��cJ�x�	��ے/z{_��*3�����g�:g������2�5o��ln� S��_ܳ�]���j$�h7֖JG|&fuD����_p�ş��_�lv����֟l�X�꒤�bN>�8Ju<9茦�c������.��*���{��@��U�Ky��NH���ڊ�yC��)x��
K5���!3uߟ��:��Մ[�d��cv�Qs�9p�b^ �cbT�̯�Г-Θ��`���9-��%A���:-�h�K�����!3�,\�#�K�<Gl�ۮ��sr9^�z&�\� �}��SV4�T�뚐���A)�ׂ�ʪ� �?Ϛ������ �� ��hk=��k��́AN��컬*��m����/Q�~ޤ(A=�*���5�x7QX*�1� �;�>D~�C�P>��[
�/?"ƫ�����Q�I�m=�B*Ht�Uw'�3�Q���ޑ�ՁKG C�խ	�i`�$~jh��S{�!/YR�G�+�A{�	�1X�5���W�p����3��Fe1"p�gs�ܬ��)zϭ�s:�B���F�vsU<�uuC��LǇ�*Q6{9v�t����[A�����naR O�q���O�"z�S�6���J,O ���� W<������j���K}}�2�{�}���P�� �w�/�H�\:ˠ�r?���h�"��@=������>��^Iٹs�e�����Y���-M�H�p�0\V�N���U�f;�����)�&3](�ع�����K<m8P|3�U��f����S���ܸti��)�R������~�\��X^-��\�i�9
A�oZ"��!�	��_|�f���E���������v�C*�	�C��ל�.]�D\aŔ2�^���/���e�� ��G������a���Ҁ;�Nj�H{EtC�ֹ_��=��es�?l�ʬ�������� �?m�N��luD���9��b��hۆ���⛹�B�&ѽ1uT��"P`0�DA�����n��OH�>q�$��t\}/���[�e� ��PZ�����������q��,R/��#�3d+�ɩ8:=�5�04�3HNP_E��n7l�k����;- �����Y�l��j�D����}[��r�|�ոg4��"?���L��\~��_!X�̂	��@y���pB��8kmp���E�C��j�Yf�%PrpA2���9���E�	���B���&������w�&{f傒�]�",��r�.�d�;��æ�<����y#У��r�o��h�x�a�Q8�%�{0c� +�\u�E������ߣh������3��@xx�l��Ǳ?hho:� �{:t�G�Ti�gl�c�y'M��}q*ۚ��
c��^fr9.��yV��IXS�E�Ep �.y�(i1]|0��T[ǵ7�d���娎U��(�*�G9z�$<MP_��@��z�W;�{.[�6������}[tk��.�]�F�c�$�Q<M�A�l+G�&�T��w�+3��!V��	��L�G�9p�,4����9��U�Sb�;�0�ښ �U�	�N�����j�>���&��gc�[��9?�-�%�v���lr�;�$��lC�˫��$�|�BK��<v���|%CR��������pV�1HA"V��W�[����f�����C��C/���3�3s�V2���>-T�rm��]I���̌M�?�EoD+��Kx2�HCg�0����VQ��n�>R �<,�J�@,�[g8a�g�R�x*L=p�n֙{�׸*ځ��� %���F����{꿺y&��c&��/��j����u�^�c�&h|����wKrv�G6�ۋ��8 Us1�ka��I��}|��U8�b�";�/Ƨ���| �<�F�B�Җ��J�A��.���g[;Q>._T�L4�=,���c���%dyF��8!�)|�T��4�Yx�� K:�ъ�����O����x�ϑ5�w����D�X�JE2���y蠞��������S��O��#��|C�^�o�w淨w���~��?�y(���`�=.?b��)�=:�Wj���@E�| �!�����!Ywh�߂�a��5��' (uSf����=��n�1"H<�v��Z�j��Ow��u8�I����t3���E���j�dc�R��-�D_b���B���k�:&0�"SY�`i �9XC���G@�������A�o̭��`�_L��>_�~����Z]i��gd���o����Ͱ+鈦S�/2a�Კ�![���iV�� Xo0
�wռ@�]c�k�I1�k�#�F��Ђ��X3$��p��Ne/ЫĴ渃��.��%����vx�9�@92��?JRG�<U��8��V����BÒ9���"�΁Q"����𡭎q0���%�]L���� �MT���|�;���k�ŰG��ہs�����2�$�U��z�&k�D)cZ�i@�/�"��f�����&'�{b��իӅǁ�x�Sr�)�: ��8�ŗ�߮�Y�� 4v�
z|�?Z���e:���(�Ưų�P��.G��4�9��Έ�IAV��XT�Q3�4�]b����8J秽j��r�j5��_`��U��I��l�[�kw_G���۝M�<�k��($�S<o;�:�g�})+��bǾ!*r��e��U��>�\(�NIɻ1��@��R�&�����-��Ă5���x���b=�#����)7N�8��2$��tEk���I�9�B�~&Rn��5F�@��=��2�=��=<F��]Δ����FG���Y6&%�Uf�0��S�={�4��hʽ�ŷ����S�|,�����������oP��r�%Z��^z�=���{5aי�H�u�"�hX����'[�t�W�E��w����o���B���������I'��Ԁ�]�R�Y�� ��0�l�YyS�yE�O8�ķ�s`=�	i�	�싂���R⛏����O�d���=ԇ�-Å~ y�G@��F�_�ioKS%JY_-�`H]�w�����`{$��L�gu����Z^\*�\�(�,�f��į��?Ƙ}֘����˲�}�ZF��s��z��;�6��"<��f�CP;I��7��;)��t�N��c�w�,B�b:<��q@H�C��=�Rk�ED���MF+��@ n���������5�Z�(\I�K�e��d=�ϖ&S"Cs:��Q��m/"5��� X�_c:'��ڱ��ΐ����&��RT��6���ܞZK�B	Aq{S#s<��^�������%LW��s��l%>̒޻ᖟ��/V[�N��Ѓ�P��~����Fv��}�;��c���؟ҁ� jUr�In#�#��y������{"�b����=6A�V-t/a;�q��kn�Q'hY��JI)��y�BD�R�����?�Z[	yg�U�QGz�j:�{�j��3�a�{My2�+��ȍ��k������ �X�X�x�ܝBRqH���9)~"�F����� u��4t����W�[o���=�Yq���h;j��0�G�dL�A�J�Cz�\���[�(IZ{>7�]�-��W�w^~��Ű�W
�б,�ד��R֔�X�J�(e�!�0t����nՋ��tXQ�
;��u��iN��EɰFG8���-�T���I�q�/K��J^�/\����#�Y'̲����kZ��g�*{%��(���4�)C��Ժ�^z��	�ķ$����t��
ߝ�;܉��0�ු�g�t�r�S��6= Ma}+ttHhë9h��zW�q�g)Q�>3٩� �"Z'��AB�&�h��A��!�3�ګ?�,���m�9�)zFR!�&&�j�h�����-�a�u�ɷ���#�Z�m��ۮ3��U�����T�֌���)���R�Bx�葧\�ly4�&�zB[��|�C��F�aB��2�J��P, �P9�?�+��[I��6b���y�R�|�V���2�^��G�:�c���6RQ ��\�N;���6s��w��ޔ�ˉ(�맩��6	�~��j�DÀ����g>3�N+7�Ә@�`�("����1B☆:�J̛�4�2�F���0r!S��6;���'�,VL���+�Zj�{fW��1|݂d�ۛ�H�0��C&�l��l2�9LyG���I���H�P$ǈ���r`
�e�:�Ȥظ�ʻQ�������aǡ��;��0��Y�����ƫ�!��.|��Rݔ��,�u{�d9�g�馑�K�|����wًݱp�j�s�Hֳ@y+���=��\(�t���/�����!(��BP<Cr�@��&rc��{���񡰼P����XYJ�yz��Z�s�U��q����z�y�y�$a ~�DD�?�\�T����L>��զ��2�vcQ��\s��ɪ�������8�@s�6*�(J����ɭݢjF�Dh���'v�r~�p�������H9μ��f�xs[7�1�tЈir`cr��J;K��#����7dC��3��c|�g�u����\�SÚo�0��+����+��G�����|��6���O�ܩ���uG���9���� �;tfM%��7˭��ac�p�'�Eq���u�����g�����у����^aϟ�[yY��u����vc���퀀�b��|��5[�NVn�8�(dn-h��w]���vF�v� �c�����Ȍ�u?:��$H�6���NN,���� %�] ��*�>�7�Z;`4���Cz8!P����Ɔ���
k�Xj����o����y�>-���
����Ty_\�p�9��{RF��]������P�B��$��N�˓tN�5ҽ>�vd�7�� �� ��J�H��D�@?��;Z�dgE�u^�Io>+�����A>��O�D?�_���+�S|�_�׷�� ��CВU�<��׽K�������q�s��'�c��Ug��^�ơM3�|�V^\�TS��Q�Xr=�R�����j��>~,��v�Yi�[g6+�-J���\��e'%DE�l��bV�*�j����ƥ�]��-�;d�<��UA���s}�������f�*%��].Ԗ��a�` ieG��h��y�*�S��5�_�9B|@�b5F[T��f��Jn���R_:�0*�؀'����C�3�}*�@�3��ć���}<lUNG���?Hp����[�ܵ�G-�OP�jW�s�F6Mؑc���H&����s��1��_���_�H�ء���z�P���/'3�E`łE�pE�80m�~�r�o,�3�p��o�6����M�1 ���}G���P'K �%�'%x_��7�b��tN49k�T�׾х���s~<2���
"Sޞ��J�"[m��/�(F�Qo\ܐ�XQ"��z1u���E��^���x�/��A�� .�N��K��S�Y���*$�G��. ,Q'�Ҥ��jb��(|5�Yi̩��]�W{d�����g�אe��
Ϯsr74Yk3ހQN�Tл��IN�7�8I#Zvq
r`�t��P@�0*W���,q��u�9khՙ~gOL�ܚ�ˡC��<�����y<T��i6ΐ�����FI�@����5{��+me���J2�k���;>g]Nm�-�1�zA�~Ŗ"�e�!�Q��
#:󦀏���0�R'㍑���w�<�)�I�������~C��FC�_ĥ1\�HL��-Sz2�I��G�����ˤg����F"�I������4cWlJ�e��EpP?�8�G�S��z[-�c��Y-F6l2츞0**
���M}ƛ��"����2�)�bҺ�{�&I�^`?����Q��v� a�u-V��//[uc�`���%i|=��j�b�ItB/I��� L�W
kL۝���6��	i1��헔�,k���g�<��1���^�}ɥ��՘��B5dI��҅���)�T��&A^�|>G����r Ia+c�w�����v]FC~N^�k����sl� �h��!4u�yhO�8��8|��9��]����E���
]�gb�]+��V����_���v Ψ����Ԃ��D_���L}��rIf�4��L�^���y(i�&�S>�)e���B.�Q�W8ƍ��Jo�n���i�_ij����|�ə!�$�<o_���ħ6�z���*�ڿ��lĩa�&ɵ�'n�O�=�9�2���0���� Tٹܪ��ΛƇ��Ş����XG<:%#��۸:�FJU�4/|�a��du���ڶz`�9vm����D����/Qo����/�����9^����&��p0��ȿZL�R�-NErb��Ӑ�O��B�#���Rf�Ӫ� ��c~z� �we��5�t������?]��C�k���)Fӷ��Y�A�4���ˬDN�A�`a�u���z��D�o|g��kkpr�z�u�K�1F������"��/x�}��qyaC��� ��N�V`:u��B5Bf���ZS
�+�A��[�{d<��G�2��a�F)��f�2�i��52se�m��bM/q����ʤ��?�<��+����J�w���y�Ll�Ogt�S�t���Ly��&�95�:�p�.���J���2\I��f�n�% :L��g�#Bj�X�\�q�ATq6x����@�� ���p������{���4��2͍uL�T���}�Z���#x�<i9�*9��߻,!����������I��b�heP���C.íƳ�S0&��� ���M2jb1��_��6.���� ����?[3�r㡸2���Al�-?޺���]��|�z@�5m0{Z�wM�e
8	d��DDCd#�!��,�@��N|�i�d[�AWL�)����Cv�|��f:>B'�x�l�w�c�.���я�����<i��l��Js����-o%�G���7���?���\�>-w�^��0.T|�a��$	@�fw�Ɉ��LUp`��き8�=������-�΄������D�-�c��t4I{��d��t3E^
��w�",�-����{�k���ԥ-Zh���ֲ����a��������[IM_��W)������qd�Wl/��0Of\)B�0�x�t��4*x�h�G�.[�*�#_��{��y��6"/}���kN`�؀}X �2�Y2>���,2��lEj�&r�"y�� �5{�9Q������h�������p2h*�����d7e����|+��'%�
�vZ��-��Dn�'\��'I��v
�G(�opts̆)偁0W����_��"u�[��)�єE��C���U���Ņ/�Q�_�Cq�q$����*̯�q�'9n�c�MG��"�vo�٩^6�{,(�����yv�4���%Ve�Lt�m�8����A�ڧ�5l	 ��/���WB���|�yWn�N}��N�AYq�}��s��q�P�I�M�f/Iܮ����j:`���{D->�R�H���r(�?�Q�#\=p�E�qC�-��T�26>�B}��7��AI�#qpa����8��Z5V�.�n�32]>w�st�O��Q	�.Į}�'�$Uk�}���@�KǊ�1Vu"��dÙ�a�q��T������Jw��[�gKS*��d6��?/U����%�R����n���U|6~�����bZW0b��o�z f��c�恒N�,s��R*��R�=��̙�Q�4&SKAN�Z�XJ���&��1�1�u�+H��ՄF>;��)�K������,�%�0��4\�*�2ve�`C����M����%i�.�"wrF��$i%4L�w����k��%K�~8E�?2���u�$8�	�sT-����?�f�@�<�l���ʡV�#�R���{�� �����3+ξ6�&$M�S*Z�:~��sP�]�{��Ԋ&�
�IEQa̫Rѡ}�e�ʏG����.�� �"�6G��.�`'��%aːI,A }�����"�o�(4��� ��,i���Ur��S�4_�Ӑ3�V�v��*-�B������l7�X�g�=�#�T��O�1��+��� ���9�m^�i$��>�yl��8�-%�����Ј�p[�\g��2��X�i�z�RIi�r��5�ZȎ�a�h�x��~'wj�?lG�Q��E��;Bdp��T�
φk��-�s*��O��:��v�Fe-s-�[�o�#�e���Tc�ط1e�)�*�d=�/�$٢ ;��I�u���O��2���RVR��W�_+c\��a�J�q����O8�:��XM�gL��o�X�X~x�=>|��B�Vi��=���}�bX�.[���Ci��5"WǮ�T��_)֪
�ߨמ�>��� �3�����1A;������@��U�ݢ�x�x��K�|Ev��(�K�����0�.��&���X��+1�y�`��+9���������Jp�p��>�čs����4�������|[�ʘ��I> �+]�+fp��Ǔ^���5SH�L:itwFKL�Jy7w�Ԗ�H��|�/���1����l�Tu;�i�m%�����g*p�-�ZխWu��%�p���MF8��S���l������hS-��:�Mn�����S����.�͂3u� >�����У�lN}���k�60��^�3���$>�����1��G�Wi@5��q�VBҕƒ�2�2�K�;�i�������ᄅ��&׾Y���ףU��J��#����H�/�")�<��}>���8w+�Z$�N��I���c�����t)�[pTng�Q�^��l^5��GU��P����IX�/ ��^0GNj���M��Qk& �ˑ�	�'d1�Y6�g����"��N��%��	1/c����p���l�2U��
�9U�_3�<�*VV��ctyBW�t��'�,JyÃhc��P��P53//�����M���e�u˅J�X��ͧ�,�Wp������=DL�O�nCR�ۧ����� MuE�V�����d��NJ0G�����v�P�1z5�G<p�S��/(da�f<�������o�	2�~d����gVN���0�x/x]Z�Wۜ��@FM�I{B=�8�ƀ�'R�L&b�s&�+��va!�Y�goH_!�q�����D�� a3����@�p�r�$����i�	�G������'{t�{l-�����B����n��eO!X0�H�Ga��n��<�L�p�Y��� ��KDw܁o���1�1o��T 2gu���	��w<�o��m�=y���хIh�x�Bujl!ExX)����*_LR�#9��S�BB%��0�
�ـ\q_.X�t���I��@@,�y��*���N��m�cfi4���((��ʪ�����|��M��O>]��Ã;[�3�W�ҩ0G� @*`�яv�ql��J�����%�
�ƒ#Mv���nr�K���������)꽈�B)D�\;���*�NB;lO�+�uG���Cibz5U'z���������7�����M�o���Y��}Gm���>�E�������3Cء��LCN@%����.g����f�_�T0,%}sƏ��9���]⡖�m�GT�
�Jg���3����R�A������xf�Z��o�֓���r��i9�ݹ�uHj��-��A��|��Ю�R�c>h�U+�2�����ǥ;�%��S���RO;���M��������7��TB�����R�{�Ȍ�_l�i�4��M@R����9���]���4r�P��Y �m�z^d�)�G�ҍS_�~����!5��t{^��!%��ۉָ�}<�W�k��1w��4n1�r���d0V���10 =	O�@k��eO��hj����~��!�U�8k D�����2�lQ�}�Б��	 ��4��E���+Q�K$� P ~�8%��M�K3�ʈ]N�����$��r	��f���O鮓4��9t7_�� �??�K�&����x�Bg����bS��׵�*P�	�~m*������O�,D��,~o�y���ZQ4{Q�!.�[x�ՓY�{�ŀ���Pݧ�u��Ye�N����v7_��(�"�Ub�%�r�|!MgӅ�怎���CI�׊�� H#���*�U�a��.OҘBJp�n�s��쩀�kŰ��Y�d0e�����7,����Y��_1rk11�%J�\*�eo�{3lPm���'�]���^�O���_h�S��&�d�����x�s.n��rb��keJ�2 ,5Ĩc:�9�\O�_�X���!+�6��'{�ɋa�{�W���yr%��HsNe�kj�747�sɟZ����B�n���8O�`����g���C��x�r�]�&�:,g���1��&�Lgmi�AP�}D���ؤ.ͭR��!%�����*�[�Zʦ��8�ԇ�"�a�'��hO�I�tdا�JR�̺�V{V,`�9���,nZ�0�0V��o�l~�S �g�ѵG�]��	��ne�M�x���9;E��UxdGb܀ �@�e���"��O��̏l��ȇ�6؃f�f�c��ysՋ��?�:�0�{�=1�^�=⥦��ِ�n3M����-Ϥ?�c��G��kU\�� V�T�"?��ޥs(��`(��́�g����%*v�Ȱ���ݒ(ä~dT`P�G�"��m�*��8F��}0[H%�G��0"�*+c��"l����sA��C�8��ʾ��!���*%CiR^ ����U�"k ��S���P j����{��Rط�n��<�E������BQt�[�nWk��nO�j��B�wg#���MFh�<�2�o	��5�����J&(�	�g�X������ �!F�heƭA�fB�*:��e���R�c���>�|�4�����3@�w�M⯛��?J�+Y<���(�o��h"R17k�Y��a͂��s�z��xǘ)�lQ/
�Qʝ1�������K��]��v��x��Tӻ~���݋�i߅��Ka����1�5W��J�y�����j��x&jw�q,��j"Я��cJ�2 ��K'��.5}H�%3�&x��Eޔ(J��%Eĭ���*��mP�����}D
W������.rI��dV�#�s���[yIu�t+ ن-"��Ms�,���5�;-έL�9� ����6Ѻ,
;׹~wl�����ܬ�LC<���KL_�<z��Q����О��N`)O�����m_|��I�E(�O����l{V�:C���^#���=��È�i�!�U�|5S��cm�CLщ��\	z;PDE�5=݃Ykk��Z�uZ�����Vǫ) ���J�\ㅴ�A,9z��a�o[��kQ7)���tr�h�Z�>{�O�Q��Z��Vb+z<�Ƒ}:����vb��0m?����*"� �R}�ΐ7�rt[.R^hp�b�Cԁ�j�H"]���nF/lN"�=�k�hW_��'0I�ӱ�B5(��=N��G�Cek�@��yL���z!��)� 
�}G �6VG9Ʃ�.��Y�"��K���:ih��|M��7�T�8���s
���Z#[W�G;>q�����l�G���~�����4%iGktl�"�r��5TF�X�h�WJ^ʥ��)��HV�Z��%T���q���CzGݍ�-�]h�"rq�XD�b�[V(?���-�I����A�c-��(U/���D5t���(��'k	Ϛ_�<���&z���.�nN�-�p�a������ǍA�l|�,���D�uu�� @�y{7= �V�N%����=��JO{ B��� m�w7M0"���~��x�x�׎z8\�=�m!��N'����)X�Cߓ�b���w�S"��*0/d�v��)C
%G���x|��%��삌�OX����jp����`��CvF�.�)B�H��~Z���zkJ�zm��r��5�^{�h�F���D�rԗ��\'8Z�7^��M�]Kqgj͟
B�ŝG@o�[4���E�� �rΞ�|��㒮m�dļd|��!v`z�CVr�d�>>�ᳫ󤴱�T��X��������8$.��/.=+	��h6{9U�&/�3��kE,mh5�[4(�Sp�O�B	kAF�q��a;��Y��Xu]��tR��|G���U:Q���{��M��$�C���	\������W1��C�C�H���ʹ6
ď��2��s��`Bv��4&#M�B�([_��ǅ��F�q5�Y���
o��3�k�p����uIkT\�A^Qt�,��I��l�pW�g�숮�W�I]"��,;���^q!��	lW`���IL-�(����
(}˰@�������zG��! �D�}q[����'h/bG8�k����d����A/s�˯<i���^�R��|)"� ���9L�+H��!�N/�S���Ţ�Ѱ"�Q/��$Tf	r�d�����X�ۧa��ﷺ *�9�#5�����6u���ߓ}p^�Ȋ�c�7X��Q�ə3�̇��xz��0��D� ��墋�Y���yr��ϵ@����u�T�M%R�a0�Y�ނ�����H�Z�[U��o����FO?��-��Kc�1��V�����f��g��|k��%�m����C�
�F�҂ƻ���9�o�yw�@�W��D��2�b��AߥQ�K]ѥ�;�
�E�6"6?�Or��U?�B�
�d�@��3�-���ff��Z(ýg�j�q�� ��Ɉne�LPh�D��S���6/k���CG�Ru}�x�X'�e�k9�tq�	��$?�y�sA��Wܑd2�&`y���_͍���XFU���B����]�N����=�[�hK�yP�kC,�Zkes�8w�C�4��CK���~
���1o�u�v>�f��O"�8p�,/�m"y�^���{`5��S�򷥷�:"�@� ���g�#v����B�
�V�0� Ƽ��5e���)�KR���c�| �v��6~4(zv��ۦ+�i�)�[i�[G�}����c����N�?�z���6�����F�D�v^��y��&��ߞ���Fw�����L��fN����u��bj�I'�m&}@���A���I�I��@c�N�#���fJ8��BB���8Z���a��<���������MlF�g��c蓇0	���R%
૶p}[�	�8����mb*Fo��T)DS����9E�cCV+�hu2ZX����?�7}��V���QGq����BE?���KZQ(q^7�O	�Iq�
�KYR�2I'��C��,�സ���� �H2���>4�s�'�?�ܕ��f���e�^��||	:��=q�e7�6�bz�]=3�+zL 7��~> :�[/,����TP���R�&����Tk:% ^ E�Δ�@�C����q��:e��n�@[���(���e�iy�B�}j,�_ �kV��|�f�������+�����O2��'�ޞߢ,�꿭D����J�����倄N��[�`�Uk��G�qMՃ���b"L�ݡ��)�_ެ} K/K��֯G-�Hz�F��cqx�MrV�}�R���Ra�C:#�ge���b����NX��Q�tQQ��#�z-��8��ݱ܍�u���;�H�o�))ЭE}S*��V�<Tb�o�u�����ª���T�Wc����/�|="�_^��5g �����>i�ܮ�9u�z�AYR��&��Ʌ.گ/^P�f�g�[�x�C��` �'���,۠��XZq���'p�35e3�K�o�64���Ԙ�?���VhP��%`24D@����|��������m~3㓡&	t��z&��4�_1_ڐ��T4���%��W��E葹�Py�^�?���.�)M�ƴ񴧳��a��U<%:k	\�|�b����^��[��>#�.`�<�:��� �/�=��#���e8�u|ao9��Q�q�6P`�`�A�~����_��b�ֲV-p܅��40`A�΃ȓ���bu�)
��٨Ӽ��>�v^�Z�6J��$^��22�
�����yb�U�c��3K��}��L�����雂��q�j.����#�?��B,�O�b�(`����ĩ�yɡ��rf��:�GB�`m�N��_�5�:5�Bָ�5i�Y���tc6���j�f��8dTAI��(;r��.���H�`��aozwx6reΚ�/t�vj��#�����g�E��"y�Xa�1�׫�,-&I���Ѫ�g�+�o�w��C���r��,�%����Pl�l+�%�Ց;9�*zA9�nc}	�=#�2��T��5z˓���<����������?���β r��aK۲B��筏�:��i�E)#i��������qa�ab���qX1�!A�@~�WS��k�����l	�K"��M�{@��'���^�Lr0�$�����,7$����D��{��@ӂf�xa,"Z4}	s���^Yd4��>�vA�S,��k���v6F��<7�����[�(���w�2�'���R���)^�K�%2�%�>�șB�����p�\�v�2��'�Cw�K��p�^���c�qԆ�U�`����*Y�d�`u����/� P���"�� 9��)G��I���*�Q����f��Xx��r������ɾ�wՋb�oYV	���7�߈��f'q��
�G^��(���E�R�R���7�1��;���-] �����E^SS!N05��'d&~!�#�YF���J��G �du4���c u��x�J�JN���n�R�mŇ��l�8v���s�lf��g,(!`�,�5`��=�Z!]�X�Ϝ-��}:��a]f~TBi��[0�2���K�㪖q�'KH5��W� ��Õ��dq�)���-�j�$l7{L_�?n��7,3*�XT?���ߗ��m(�ێ�$�N��}?�gd�;l�9*�GNj��x�:�#��e qR!�I����ƇS9�g�N��_J�_�%�H8$
W ��tx�[���֋Ž�Š��D�oV�Q��t�5�7�I�����7rHv
���&I�Aзh��L���E���B����BZ�B�1�9�p�9��i���SM6��~V�3���n�4��.�Ff��&���|Q����(�4���N�:��[��u�\�Ƹ''�Sp
l����*(�ZΈ~�3���9�!�U7RH�~���:8^�&�=+��@����4n�t�����BP�ɻ�\��i��!t��;�>/D��R���l��%�ȟ�gDA�T(�6]rQw��sv�k���1�FG��q���Z{������%!�7��<|9W����5ĭp"!5��˹�I���.��e��&�$Y-�r!!|{z�f���*"��CUNΊS����ّ���x��QKT������'���ÿw�*�ͣd6�兌�{����Rn-�&�����$&�7���uai���?ؼ�k�a{���V�ԕ3zT&�:&�X�HH�M�w:���x�ݙ��{�mo��āyp�^2�����
�*ƒ�n�cLG/�Ӹ�Dtz����>Jy�O�i4G��+"�+��ZK�F_����6G�/�����yT���Z@'.�pf)lt��tx��4�_y=�dY{�[�l�\<�1!���\����'�"i�p~ÏjJB�8	��gՐ;b���Q6/+k�N���
h��$�O��=oj�Ͷ�{�c4�{��@yS�R��&-ac �qL�y�)����x��:�$��6g�Pt�1G�jہ�a-G�U3�&a��縙uif����$��¨A���)Z�efލ�f�~ጏ������G1Z�C�����}LJ%����bd��F�̧T�{v�ۃ r2����^C�/�|	�	����Eޣ)�����:r���u�����cJ�E�ܯ����6�>96���-���j�&'��$M���U1R=Bߊ���dN�m�cs����ѡ���޻�?�j��g�'��qh��4ӎ@��-^���S#�ZJ�7������Q�9�cγy��KK���%A:���lzD��#:���آ�Z���1�s�%nUi��(B��� �/�f�Fc���6i��H�/�/ۈL���+X�ph�n�4�P��t&��+R��r2,#)N���9�z���pH�=F"���lT/��4_�#�H��FD�����@l������+��� ٮak�,$b�s�<�$R��USo.�H5�9尭#�ѷ�ۡ�x"P���mP��-`^&��#�����6~-�>����\;�V�5=K��,|*,5x�>��fqf�prb���ul�[�>�����Y���^���w��7�@��T�5����-/<���y�|Q��a~����,K���x1��6T\�e�=�o���o'µ�X��p�u���#ys5d��d*��k	��PҠ�),�����y,��z�=i<�B�{�������(R���N�ko�Eb���Ph�H���3�7&ulB�j���G`�qD�@|�֐���2�T#Uq���xt���=<1kUY��F�j �+�6�yb���:h�0n|������l^l���`�m�-���z#��ќ��]O�Y�Y8�����#�]���dy��)�޸B\�wÚ��w�@.��S?�z4�X����K����M��˓H���*�B�S���^�p�p��I"��,�:qy����"����P/��xu:L��þ���I���k�s6�-I/(�np��.���u|�x�x>g�e����h��[�|~�F�pl$w��-;�l`�a���)�����P��'g'���ۍ�a���Hz0 ��/�a��>�;ɨc��pr#Z�j��"�l�M�	K�v���+�'n(@�o�k�l�6��o�h?�@hb�6D�2�J�U	��&p_/���h�3��I�h�"�v���B�=ꏆD�ZU��M1��zЕ��CV�����^B�>ì���|H#��4؞�$va��k}�6�	Ly�� 	���6�+I�}�����A�%8Ǽ,��Vw9A`�_�)H���E�
����p��[��+aU��++l�{�{Fx�'�~�.�H5��'�cZ��#�4��]��c�1V^K.":���CL>����
p���Ӗ	��/�:Y�R��`jX�C��l�)ӔOsKj'Cפ@�����0��Y/y��愼�>��M�X�X���ʔ��3��л�w��ǻ-��ƐS���{6���UmK��J"�|�T�K}���ڛ?0>��>�eRDi Ν�|{b�^uk��0�O"1Y�<����P�,K�#�z+y<�-������, 瓕Kn+��d^8�<���K&������K}b��'������o�yHl���s ��}D�5u��׽�71��N�w`ʼ�-.,�7���)Va�x#�oyb2_;�r�z�'��������Y8^~f�u�(�б�0Z��٬��2v=�7m�&Z?��;����`[t��\�t�ӟFbs�k.���nz{v}F_Q�-1b�&��3���n�`
�����!�P47�x�^6S�P��m�đ��o��N�<���=��<�=h�cU|���-Z��z��%h�}�犘o(���h4/@��3�\��#�����=��c�<@!�\8~	s�P���3|�z�ܻ��v2�mJ}'�L�q+�������"<aQ� ��ω�Al��-���7�0/�w2���ح��q)C���������V�\�x�[��Ƙ���ߺ�
���Y@1SH�,?-���s����Y�蓣AsP�ˊYͭC�Sd�hc���©�S-e���g�h�o�8��"�b��P8����_w�$5��h����B��ă�[w@��7/O�R�u#���o]�����&�jI7;����nO(�Hx�b�&9nC�x>��~`���%��ŷR�P���-�`�������\Pf�bl�҅t�:����J���)���kc�l�&��R>c'�I�7���_u8�k|��F���n�fS��f��v������穢����C���<;�WL������ډ�^�����Tf�m�~^��K�Kdf��v�'tP���;�7�l(~�_����V�5Dܮ��nNZ��}�[�٧�� �	��;u?�3�@%[���=a�J��	/�N�MH�;m����j���ok)�n�� H�b4��'!��;=Fq��qJ��i}{ӎ��/o��u�0�a��DЦ���}9
؃v�$�V!�sYܱ핱RgK�+�dr�7�~�R#R1ԝҬ@��ǆ�㚌?�n�Y�.�
�W[�O�c��2.a���E�M�Ut@���,����
I߱ @*W3��@�0.��/ZA��h|�DV��y;�WC�#>��^b��i7ļ�;�C���ެ́�8%�K���L_� �{E��zn���mf
A9ڀ�YeK�F�J{1	S���k�̓2T��Ɍ�x������0MFngy��\T�������aY�啇�N!?�<������!Di��ǩ�����X봱�Xf��z)i5�[�j�_�`:�k)c�1Pt������ �ݦ)>�ۢ?�F��]��Ѽiƀ:�8m@��D�+8!�ϣ�!�u�~!ppj�B�/]����/���i,�f����U0�]7u��ya�氛�:-�^I�H:���S���r�&)����{uO���%�]�`��sBO�7��3�N!3��`;B~�����$��~��R���Y}s˶F����M����C�w�Z�i�?�ح���`�j�2z��Y�1Ŋn���g���*�*�8աXWǘ���9���lY�<C`,�|�u����U��=�j�k�Մ1���d���ɺTP��.%b{�t�o_SM�`C:�B��5���5�����PXߒ�5�v������f'��%�T'�(P"Ö-{lADM�]���ۿ��tmD��NUm��R�&ϻ>߬�a0��gi2h��������(.���:��(a5G�33(qPξ����1��N�f�w��Y28�+�y�~J#fc1ߍ�CY]c�h�3��t�4�=��vK��Dp�Q��R��FHn8���q%je#d؁]Je"���O��C��i�SSg��>S�TtM=�'0��J����W��L�W)�e��Ȥ��J�5�������a��Z��NW�vG�R�C�2	�[;e��*�N�!���ԑf���s���[��,�=��f���# �{��l�o���&2(���%^k������k[�J���p}�>�Sg:�'�풥7�U<T�c�M��B)����	3�{���N���`�.	��t��7��p�6j�܄ q*,�C���6����eǋ�^���!���8�AFpT,O�B��үԖ�SP������٬C�y�$�V{ $"Q<�ZFA!w�ԑ84�{v�Nߣ3�r��[�Б��(n�N"v2:3��_%ĺ]��e�(F�5GK)��7�%�2���~E������C�S�UG����ȱQqL��w���H߾��{D�C!�R0�0,eM�b2͛��I�=�ŧ\\��ڄ�A�>[�����Kߝtǀ��T�3}$�_b$:)��P�����ϼ~�5Ⰾ�
��T+x��)d�P]V�r�2;�P�S����p�GRJ�.�f��ާd#���b֫c-�w�w����S3�Y��H�6Ӛ+屯ګ�6-��(����\��A�	�j"����C���A;lWZv�ҸskoLgY��s`zL��ÂxM�.��fi�Ā`�7�3�B�j�/�ٷV��9�qߨ��Q+�Jw~A��yL�o9�9*`�!D"����Dn�>����HpN�@&>�[��Vӭ[El�_���צ� �Z�W��m�� ���A$�@o���x�FF:��7���q�z��.l��1���v}'?C�������%�����h�l�d�y,{(�2�u���	8�{h�k�����>m�f&n�(jh��ڤh[%�pй�������{���!��	��(�/�PY�g1ԠS"�"p�Tf�!B�5��.��8���m����"8�	�"pd�	���&C_�:3I�f=��ょ�{���>�b$ъ@	�t
-H�R�To�q?y&8�����U�6]�Cn��5_
�cgKLQKԮ�U�l���xY�V��9�6Y�KG`�1(�����?�rĐ�OG ��?|+vИ��j$�1��Ѓin�`�^��D����&Zvԓ��4��a���Ƕ3?��E�R`0�e9TR��%�P��W��FI��K|wIG��uf�������Hq�����ڹ���}���ʑ�
�1\�R�uJ�\ )Y@�p���a��|�	;�?IR�w��d8�cˤʬ6� ������G��PVn󰕈���|��9s�9�n��=�!��o/�5T�ŗ�"�\v�3�FN��ml&�Z!X���]i2��{7ӵ-���0%�mPm���z�s�h�6�kّ=�e`'=��.���m��'oYކ9�J>!�f���ރ�` ��P��ԏ���������K�l�>o���BI�.��t��L_P������]���8��Z�ɴl��{5���2����Ie!�(�y�n����^	�e#37�K�ڻ�z���m�Jl AԁYC���R	n����c����Y����� ��*EF%Wƀ�
��s��rn2"O+��J�^L���^�`KaTK�h����H��Y��T�	�7i��c߶翦�
�� `�XD���y^�<ث-l�햹DV$ì}�B�=�'�JI2��y'�OȠ�A�Vkũz[�%��leb�X����&3@XS�)q D��������-���<���O���V`�+�N��,��/!�~j��8���lUy��x���X%]z��R����4�)��j�`Z~�Z�ҏYrtG5kQ '��>c�+��Tg���o�t�}@�f�]�2�z><���(�EU�q"n�,�~eʧ�8��L�
�SB��m��+�[91Q,M�V���Ez^<��7�_r�J��X�}B�
�
��	��2n�P�'���V�ve�_��O�Ȩ�T���\�6?;]Tݍ��I�f��R2K�,��`,<s(t�Dd�
U��Эm���I~C�<�� K�$_E4�l����=�E���E�S�|�'�Bل�*�������fu1�RRv�޾D-��>`�QQ�K�E�� (�qv��4� �w� �":~o<��+S_�/���ӱz��W<�+c�kN�I̩����S��	M����.k�KPJ#����?2ݳ��V��q躤��w���>��A52\�: ����(9@�0V�v�� ���y|��92��=�oX����Nj,����)�6��Q�<�X_1�p �H?t��X_@A<��Jj{!�JY#� q�c)<����t�lĝh���&Cю'͜����~�g�j�*���/9ߤ^Į��_��:�v�F�O3+��j����Gy>���zi����
c��G�s}�hUFy�u��\7�{m�BQ�Ն`+�)8�$!�)(�]܃�}A�4��RdLe�e]+E���2�~=�<�]�5C7�`��o:��`<���5��3|,X`@n�_Gk<��5\��J��nsg݁h�\���KB���c�V�F0���?�M2��zIoO2x͸���ߏGmU"r��u���u,�姘 �Ih���D~1i�Z^�e�<h�����s>@��
E/.䢧��\��o�mc_%S4|�Z�5�j���wy���i���`�\����ޘ��Οh���N� ��*����4���;x�jo�k=d����!��'�C�I�]��x���C1�v)����ʔ�#5��5|"T D���<�P��)RV��J���	��;.HD�W'�C���3F'�w���!�� (�1Mg%VA�*��	��󥦵��E��Q>�0)�9�{���C�J�*��7�~���C,ǞUm����h��������B��JV�@/cX"��
udBH��}��]X'b��
�������`T�qɝ��2e�Fb���h����U-�R�$314��Y;��IU(���҆N�~�����<���k��4Lm���ԏ՚�'f���T�f:H1q�\�?k���I~pc8e&�K���,����BD�o�f	 ��>��4����q��}�xg�(�4s>˧���VMcR�Y�˔=�x̀����r� u��j�u@`]���B��%O��\ow���B�88ɚ�(RUJ�jc}��_�IE���qP)��^���{��%ND�\��5�FZג�H��֛�@�Z�kio�Dɒ�C���H���������;�x��vp�
��QF>��%~d
E�wS�G�q���6�|�_�Sd zԢ]M�
 5A���x+��哆���4��5�1�jO��o��T��=�O-��M�#&�x�q�cǩ�R@$��u"��=��BΚ�b��ʞ	�O� $��2��.+Pv�9L��2���Ⱦݦ:�^p�4"�4���{=��y�{���>�X�5� TʢoG��XT&�-0)s���.G�-����fbFm^�N����l�z
�z|�xm�C[��Б]��'vSA�R��Ԉt�C�}��P�h=��y?���'�4nd������j����P�����/�iZDx��&/����(H��8h��Q��A
�X��e��[�@�
J8���ؒ�L8���n���T'����9S+�l���R�ټ\Q�Fۮ��0�
���G��/�}���(2b���.x3�#���t&���=����?��#1i�1
!&g�t9�5A����Ͱ9r��~ߛ���z�z��//��I! ��*�S>��F&��g]��Y��V�M���[���ͥ�Fp�WN�gD�"�<ɜ�`k�2�S�.�Y�s9p>P!�.΄c��}X��{=v�����`��Et�3��ȧ�h�
 �CA&H���&���[�h�I��ZN���?��z؆�5�[�,�(��3�F�a�8`3�?࠽Tj-O�� \��4cܴ1W��
|� 	���NY9�ͼ�]��؟�-z'\�5�j��<m���hF�o0��$����@�e����f�"�r��wXxo�A�\�~���x��ܯ�*Ket~{�	?�5%����R��uh��q4F��iqd�@�ףT�Z���:�+��)�m*Zꦙo�⥔��Z��l��?�|�a>{��Pl�_��e	P<T�W��(�(.����0~"~��GQ0GDl[[���z���'�C{��u��L����T3�����2��4�g��-��|A�W���
3��z���܍�3tm�s[����!��o�m��g����&V�I��^���w��~Q��ʲ���汤wY�I�^M�!�7��m��0K/PZ�rI�����@�
�=�ƔW���->��W�:j�FO�[ַ��PTД���DB7�2t�}�脡2�-CZ��cl<2����Թ�#.·�E��TϤ�|�[�ͧ�ڛ�ѸA2;0��/ű|�{��mQ��㩯-0����Fw��H�M�7zUf'�L��
_�LK�w������[fS/�Q�ڲ���a��h�N_N�� 3���^6�����7��ߣ~xi����F����%W�9	�/47���
Z��i�TjS�8b٧�ԟ7f%ޖ�dBh���@߄ut��^D�0A�"��i!�~u��\s�`C����a�'Zq�����K�bkA����U�n��ҹ����	A�K��S�#���F�e�Ӳ���3����L�x 1�?�&^�Z�0x��sX�ꯉ�(��!��T��FD7��D�S�9��$l��'��Ƞ�S�S��)m���9a�S l�t�w�U�Xk���<��#��A�g|�0����q"�簊�\s�<E�qqv�fP��+���>W��V�,E=��%�~���<�����0o�O -�3W!��+�	����j�*�ga��j,�rf�5�s��C|p�ڈ
S̐gPǹω@�d(�,�����-%�����B:��TR�Ym��
^�碍�8H�TI�	��A��K�*Փ�G��5�����fh���Cu�A�kp��K�ћ/`v[w��S`<
�����9ԏ��ؤ����T��a�%Q��^�U:Q��W�2I� �9+�`�<F�������j�#*P�o�j�hvf�7��<���d�X��/����P�o�҄��	i�Bez�*H0���V�<t�\A�S	�͔@���9}��\����R-p��j�@T���/�l� �G��ʝ�n�|'s�bc���q �R?j��[1er`H��is��v�>Lm�?�9�@` �V�	�6	�t�;=�8ZcK��EuHw�@�S�=��c�W>����(
�T_�����޴�
��p=��2�~{�4fYU��An�������~����p�p��brW�z����Qݗ�CQ�H�F_�v�EPD���M:������c����t�P����ލ霛��N��r�^�9|�7�~����i�i�x�x�Ε%he~��Y[�=����<ԗ@�O
1QR��/dS֦DLW��i��x	�D������!ȿ��_8�(�Vh���6�9����Ja�4F��xà��x��)�zIs��+�m^9�����0Jq�z��A�M��j\sq�W����mo���i{�`����D@hܭ:�ɶ�J�b(�j��!�^�k0�x`"�UKб��G�{8�@��	��up��6�F�I� f�e�q �������~Ằ(���c��	�s�X�%�)�,�o��&�pď&������:8�-�ݺ���s7�9����3���3���mJt3j�hN�a#���oJ^�\u�~���mM�2���Y��ǖt87���C��g�?�@��h��4��;�h�݉r�ey7D�߳�H4��h��wV�g!����"�>�=���(W��
��G)"=3��8I	�ձjb#.7�jN��D�Wo�Ra� "��Ύo�����8�h22��p�.���FP9I�AF<0��Ky�;x[	,���dU�5<��	PNi���JJq�v���� ��Hn�h�k�)1�)��s$	�kڞU��*�BAm=���O�᪕��?�|�@!���A�xE#|_����K�<�q�Ǒ%�5�ډs���&Z���ut��3�ؽt�W�u�)�{E����@YD����@�b{ ���g��Ҝ�l(�����d�<�k��_d</�5<�&Y(�[D��@�6���9�CG�7JZ�*q?B�1���a*2u�@!6 d���/��D���|O�L�IC��VM�����ܙ�{:�8͐"�Ղv9�����Y�D�>�a�p�m��������;� � �k�]��+L�i��G�pђ�|���E�+��j�*�bH�{��g?��W26�}��W�n���@:���Wy��M2�Qɜ��nS3� �h��F�~\(�a���P#�v;cl�v��q0VZuC�A<��_\���\����G��� �K���sG.zs�bn �T�d����ۉ٬Z3�ki���L���N
L�^i�mĩ#�#�$;l��(��G�W/e��3v�3^fW'⻍f��!ᆐh��Cr||�2�����(#Z�C��cr��Xy˴����� ��ip��=�<>�?@�1<7��U=��*��w��c����u�sK
�7�਽y-���vx�2��	���+ q���,�w��C*�VLbk��T��`�H助\�'$�B����y��8h��4?���&�e����F����~��'�'�t��Z1E�r��W��uB�����K���z��yh�+Wq{��4l_����`��\@}`Ȍ��Z�����wH�����'+�DE�	6��]Ik?� VD^i�G�]Ư��O�gKFE��ϸ4:(�^�OzD#�,ܞ"�z>��`�_T� �!�����9���ޢ�Iﻪ��uΝVPI[�HV�G�3)h���A��@�����ԕo��;̣���̞U�~��
����fQ}�ib�����(�	�u�����+��0����g��"g5�
w�͵�A\T?��Ա�����x�{+&iq^�u� {I���h��i�%Ֆ�q���m4�g"�,X�A}Q�:O�4�Y�/���4��[��_�+V(S{uđ����� ��`!\����J��"��'s��t�a�����~��|��) �����N3i�S�T˥%�b��a�>���G��bz.(�~$F�ת�g+L�3�Y2���h����s�VaG&)���<�$��7�FS�K�{��E|�Q��N�f,l��ɩa#(8�b�E�b�]949���q}��Q�`f��sv��ȝ%�+m�A9c��@&ӭ�y����ݒ�(���|��ݦ������	���D���K�
�Rr_:��g���)~�Bdw�n}ӀN$*��=�,�ۻ����7{���Ļ9�b�4�:�}9��#�g�}K��t�F�V�/�M#H�J�r0it���a)4�7㠮1:-t������A�F�f�ω��ȚD�.��d��PJ�CpB�����G���ӎ�+(� �˂ς,1<��~��$�Љ�B:�y�*�^ښ"�ͺJ�t�X	�w�s�3�4u�����@��q��\���<9���й�f��zh;�dx;n�cY���vpO��:2���Ǉ�E��f�4 X�B��?"~}M6ہ������+�v�F�[���H�#�f��ȟU��6��>�C��YB��kIV��絧�2z�o�����)��v}�-�D��M(�@��o���%;����[��2���e�ݽ���9^Lz;��;[ \o6bB����1�?4���uuq%�@F6�����ΰ��EAR-5@��pf�*bW��*���M�CD��[Z��]���ef����:O��l���1E��C-���Wf��`	�6�93u���F�|9�z&�|�ߪ4��c��%bˬFӼK@T14m��)���Bc���86Ɗ)�����s�F+���m��ɋf#O2[rL�G�Q��������=�|N@�� ��Ȃ\����?���rR�5-I�'h�6/���m��s��Q&�d�F�}t�S��mw��д��W�2r���r���N�= ��4Ⲇ���&�	�]D������۶�h<�p�A|6u�������}+��'#�\շ����I8p��;��P!���7~�uȗ�፮�{�5Sw/Ɵj �+��˓~��Ҭ�U�l收7H��r����#z�]��+�J1�^(���1͆_��Uڑ�tGi]q������Z�'�c��uuu��Y�D�?5Ɠf�b7,Y�<p�ۦ[����d�&���/��GY7O|�͓���9Y�P��`;�o��j�J�W)�X�AZ��ʽ�]�]��F���u���:�.������I<��^�	��l��aP�l�k����V�~}᠟9����r�^�P�� ,rO6:q���bW�Ҍ�4,Ɣ+'~�='��J��6�Yv�n{Mx6�;FR�i��6�3F{s�ձZ�H<���>����'��i�9֔%�\����"9���y�=���i�.��u�u�m]�D�%���uIE�5�E��!j�&����oH/�4zX�T0�Ʉ��=��u��Ku��@��q�\䫪S��mЅ�-���? ����5�g�38����ψY?���=��R-����$t�]	���?�A�qE��)��l�	��Q��f��N�;������Rd~As���v��s!������A��{{ݛ�����r�����0-�r��� a-؎���\��$(�;MV���i"�|$#
;�
37�&��l:L��.FGi'`T�U�{ឱwD�	G�m��0h����SvTm��|�����9�o>�����e�W�,�{��A��N�?�Mw��b�5�$�E����VI�끭d�s�3@�������Z�2<�E�	}H�(�F�rE6���!�f��?��vG�~G��Hu���_j�f�/�N"wL��,'��B`p��6u���aޑW2Dg��8��r�<�� �$����rɾB'{�gm�4Y��p����9�=��Z
�� �s$4�uS?̀�}�u�e �:�\�^v�rc��Zvc.����]ղa)�fk�d� \ޥ�;���	�w;��bզ����/�z l��EE��53�>��9���ڒb�&[��v=En��63O�:��!@�^9t�j��$O�@�r���3�#y�L�&y Ga��^�y���dV��nx�Is�&0۵ �D7��2'W+�{l���f�{��׮������(�����v:���B�������`��lc`T�@�X]�.@�;;�p:@?T&.��k��z�ENQ��FDj?��	RD,j ��Q�3u�FtBo>S�3q��	�F��©H/�~6qR�L��;9m����~���04[��ތ�RM���Fߞ�1\,��� ���े�3�jS����h_CC����G��W�=�x�X��k1"�������C� V�/g�<��X`���L�H#ـ�[���f�jI��$�~�� �=A�I�Wy$�~-��� 㔶����4��\�ݻ��Q]�ƫf��2��w�#Mm,��hNα��U3|L�����,�"�y��״x�}��ǏG1�ݧ�R�����j�����qu\�o4�G@�Q�"�!��\᧝iV��/x�2"��	�S|b��.:Ͳ��AkV;Q��ɪ����l��,���(^Yq�P��d�����yw��5L���~�Y'^vߴ�m��z�ծ1%!��s
����󼚳��y�^�����F��Gt$Y�T�����0%���ZP������r(��ﮁ��� �v1��q��w��H�u���b���e����G�O-&y6C�ЕG�E';�;���7*5bD�q��(�Z���t}᫝ϗ_ �:������3�,�p�@�d�˅J��B�u^2N�\	��w�#<��I�0�/�
�LҘ��8}X��gN�UM�:���2u�����
��� ,�04�QTu-/ʗ�@��Xj,]gv�����J�1O ��P���B��G֩�����J��<G���Uu,��#j�^��N-�a�9,Q/��m�U:Ď�������T��}���N����|�/>��BUv@Z﬙(�@t}��mNҏ��x�p��R��U�Ǒ�:[�~�v�������Z�dk�b�vȸ�@��h�餪9�� ��t;�ĉpI�qV�{s���������/��,&�0��y���8�����舍B�v*	�Y�c� ����ݢ�-�\�B��2��x~�����2j>�g�a���a�'V����Áv�|�rG5K�JG�`�V%�.����[q��\��wc8�s��ᡗ�-~���E�j�� ����ږ��멯<�0�vy����Ι�#sA��i��� �'p��h:/���]j��JUn��1���\�V=���Rde�y7)6�� :`_m]*�꾄`��xC�c�\��W�e09f�F�~��8;���Z4��C�U<���~u�%�1��̤\X���y����e��������p�S�lwʪ�-�ULy|�%+b�zHuc��G�%|��r��sUCv�$kz/�輍$ьрAdZ�A�~�ee����Bn�<,�{�?)�~�CekT��ʘ?��⌊bL����@��)��@i㳩�{�����.��r]ᐑu֢�!�=�:��]uyǺ�����L�DM<w��2Vy���v��IxV#���x��э=gZD����y��jd�f���q�Zy3��B!+�?M�����K���A��a�ق��D����Z�[���y�p	��':�Zih�������$W2} ����̧����tr#�H�? �n�ܼ""K���5� 7�
��zE\�>�W�^m;-�������2e\T���nӈ�Ò{��r~^���%y��t�����IzS�~y���O���^�w�v�"nu������ą51SlX7��.����ؚ�(���C?M�Lݿ���X=~�_g3�,���6������,McO����$N�j��VB8�m̨q�ܹ},NíxZ���S���2d��ƾ�8����#TAv��3�J
�؈��)��F\P�h���BRϷݛ�[N�y�9R�0�H>�ku�������^������KY�5M��i8���G˴#�X˞�@FP"-�Q4Mh[�ŨB�����Jl�&��L1�ݘ�8�[��f�	������ �k6���ȍJ:6�(5I@I��"��^�K�8A�f\zu��Vv�����{"E1V��=�-In1�[\�{�����.��c/��RѴ�L�q~�_C#ìo
_`E6�Ь�/���n��뗾������upk�sL)��흢|��`JL>|��p*HĔ(Eղ�%[���gEl�)�v����ע�Еw��ީ��K����XL�F�{;5߻;�l�m������yjsS[�$�Ⱦ]�Cڝ�غ��=�����U���C���`����<:~��v�as��7H���N�%0a�~9
�$�5���J��JF{	�	
��5*}�G��U�ߜ>�<m~�v"%\��	�__�_��+i��L��uL�'���[�ωZyoC�BHO�
�I�[�x�Í��B`��2��%j��]�3yO�@r��z�k����Z
K�s�AR�^�N�f�]�\醈�o�m1Y<�tl�
���r�`��{�?,���e��S@��>� �yɆ?wkC���p����o�YA�<�G�,hs�F��wc-%���.�u�"q�$�eZ|0�/G�� ��&}��UlB@��μ�r� �q�p�JV�6�Oa�N]�~�\[eԎ�&Qq��;��\ȩ���o>{ע�F�i�B�|W�C�_�<�rjG���k�rU��iy�w8��G�a�1�F��<s�����+�^;��qz�@���^^�Cg���e���b���p(;�'����%=��G�`����d��תּD*B�u�����;��˼F�Gh��W�Z�C11%�c�F�y[����P�V��S�&�\�\�fJ�'�!�\��s��LR�I�ٜb~��"��2֮���IL���RfZG��(A�|��j�a�<Rd���ؓ��䥀�����o�IC��0���%Dh��'ߺ������s�ݡC�Ma�:J�ҥA���^��[{�F��!�����!�w;Q`씀�l\���.p_F|odN��@�E d'��� &I�W�5�W��JW�e��|��a�JPc�"�i����H�\%A�i�lݔۍ�S�2��i�`�kq=ɡ���I�\x��4�E=�k����ѭ��u �
�)z�����pY���qh )y��
�YG���^��%cp��y�����}��@��F���.�؃�o&��Z��i{2.�y��m�N.n�'!���I���L���� ���� L	Wd��n\����J�Y���ȧ)�:
25���l���sy�iY�!�?R��y9>4�<�3����;�r�@�b��{�J3�^�{j�F��n'
�/��2�d�����ys�#�"@���������l#�XO�Ѭ�����$�@%����3�+π5�V���=	Q <��Y�gg�Q��`V^]�S5\0��p����ۘ6���Wφ� ���h,��R����r.�b�vFV�p^�5�'ͯ5��,j(>x�|�4vC��0|c��;M���P��2~��"�8L'P�SS����{|��]��A(�;
o3P(T�؍�E����
�'!������.�"���?3�!Ԏ@IJY���LYgJ?c�Q_.�T����s�%��e ���1�:'��~v��jZ5�=��a�)#J�z�G}�P}Ql�5������"z,A�N9IsJ���/����Nuړ�"�H�z_���u��o��XaG�,�R�O�s�e�����mzA�2�L\��8��ֻ���5�h�u�z�_ؽ �]�sF��U����ED������>���]��!kb���:��]�9��&�3`2Ұ���t�-�(��6N3� ��+��w��M����[�cw���ڲ���ҝ}�R.��$j��$*�on�&��>��F��eg���4(eרfL��>��5���9�l������;F�`�5p�;e/�7I��\k��#���Ǉ>}�zl��1Uc��ȁ�=���cT��U��S��0z�@!�d��7V
J�v�t�
����|�	�oʆ�w�k� 6Л̬DU;H��,r���K1S�7�iU�&#��Q~��f��ig52�4w�-����[Pv�u�>Wz�W�=h� �u��/"Q"nN���jc���IsS��bZl���7�eUL8<�^�o��mg(�#���d���$�e��<o��)��d�z5���?mL���-8�"�
h����مE7���)�<,7g�.��8�T�d��D��p�ETFC�ԗӨ$��
�g�嚟c����m��!�ףi0əUh÷M��4�u}�����,�!��P�0���T&Փ5,�'�n�|L�Y<�J���|,�g)�<(�m\��]z��D��݉�����c(cp���Eٵ� ��bz=���s+��{ny�8����c��y���m}��A�j���ؕl�	ۂIP�R��;1�[/�Y���ȖM� ���U�i+r(���)l[������	�7���;��VJ4H}m��m��CeF�ڢ~�2T�g����-	�����	⾢H�K�Ǚ���73�D|�h�W'��׵�-3ݯrd��l�^c������J�