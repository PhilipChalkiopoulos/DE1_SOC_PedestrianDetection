��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b����K=&no��|�g�A���>���cçс�Y�y~��5�L� ިs�4 ��ۓxd���� �9��ޗ��u�*�%QҊ�N��9��&�5����H	�=(�`�1,|lb�o�d�߀�J��"�FӦř�A{<@��!��9*��c�t]J��W�vEj���vVk8"RXK�|�=#ͪ�x�}��M�_�8��|��wX�p4hqJ���`�M~1�Ǽ�|J��G������]+"8W5P
xNCb���˛�͜ �df>�%rI�h���s]Cf7D��_+[﷜\)u��۟�x�$�!@�
�q��T�VIRq�tL͐ERڮJ�-�g�.S���O�x��h�]��ʋ�M#�r�3��O6��x�ɱ�m�ӇY��#� ���w��U�d��<�y��f�e(����\��������S�}��TH\)8���uI��O����G�f�`������?����,�`abIЋD��E�Ak@�����/�W�G5�O��[$5�� �U���m�aq��T}1��T�����E��+o}��(�9���<˾�K�g(ԟ{����
I5Q%n�F��ۂrhI�Iڳ�����)L7��+�g��4�ǽ�-���A$)��"Q_;,�7Dr�1A������8������!�>�O9����	�y1VH�3�yċ��i{5�Ɯ����9*��L�yC��s��	�r���Q�q�	9��4���}&�֪@��9[�����B�Pg]����6,�B���<m%j�`>�^7CF<��3�'���M����pF�K�[�Wx�X&����-RX�>M�D(����޴��S��ۓ�ȶ��=3֯N��o��d�Y�M��B*a0���#�z�l�r��BKl���Y"���G�����A��mZE�GzN�zϤ0��vwv�d�1�BQ3BOO{%BA\��A�ǭ�(�d�Ѫ��
�΢��U�n������[<n��1����{ú��3����'���A���,�o�qQ�L+���U��.߆��v^�5`���y��7�[�鋇���\Q�����L�$�!��i�>��{�?Y��V�TA>3��p�3d&�Y��1;��cL�;ڰ��L~s�!s���&p����;�~S�Wjv��	��J[Ĩ�E/6���'�9IS=�º�Gw�(�>;u�<�Lgj���\׏t�4��xݟ?Nҍ{�3� ս#(|"m�FA�}7R� vL_L��3�mQԈJ"��q��K���@&A4B���?�y���$8bo�
�q�(�3���8H�׼h��-�|�J�[YU"i�=�}�]�����z�Y��2�x�fY�R��\�i�m�c����c5�;z!ظg�	oZs�/�	��\4Ye�%���T���]e�� �l�23A��+���4Q7	[��z�vy#5��ފ��@�Ҷ�6���uE�b���b�\�P��5-ӵ:���u����͠�ՔX�E��ۮ���k�gS�f��݊@~�1��I�7���,j�k�����H޴��ȩl���3��a�C�:ZU��
��
���Rh��X.�����%mqD����g��O�G��S
�@
��Υj�#y�b|�"���{z�?"�Ò�p�D]SF+3���<`W��l86vr݅
wzj��USf�.���A���v��D ��߇ 	W�zp��/��U%��d�7�`~�rh�28����<�ץ��n�)��H��b�)Vd;�u�
�,X��PQ�������X�4�Ie��J2�hoN6�.3_XJ����Hl�E�A*����{I�|�WQ��C����x���U��$u�IuG��y�jJI�xQSl?Q���t��
���w�;fԓ�+Ly�^.��#S( ���ǈ+�b1$��p���:�GM�p8��x( N��*�ɮ�?ߗ����O�M��ﯳ)�\�(�D�����0&5�p'(mLz��c�W���F[��ם���@hd�Oe�]T�ߒ��-5wĪ|9��ϴ,\������P����d�,�}�������T�{Qe2�������ab	C"���fLȉ�`���Z
���]ےm���?=�c��H�\� ���B�Jz�#�G�D��}v���:租�-�=���6�	�����;�i�7��g��0J�IW�"���_�Qx�F�&���Ϲ�Ѣ"��};�:l+hF�a�8%F�@�Y����UyN��z��MRm��h��ö nKy�]CyN���C�b37[�!����t'��![����[&�F����1K۶�<�?(�C���a��,$�u����'ᘇ�~������7�u�ƌ��l�UUe�B(�L7}w F��<�W��?�h����NPh9S$pQO6uU~����#=0i���P��4;!��]4&Kğ�&�*���ۨ��pN[�n���l��~�;O���8-/,Ptv���~�� YHq�uG�����G�\|B���n��Y��U*7w_bo��aA&�b�����(����m;��|�ňP����xSR�Ţ���?�7����D>�Y,�F� � j��0��o��1Qh@e!��Ȓ0��0���OJ+
Q��A�S�"�?}ߠJ��<�m�K����)��S ~�f��	|)%3�����_:a��Y��I���|��r8�/?�7�`�7�C-��cN]�g�yb��7�A�,��5.z�>���@5�Ve��G��Ld���=��S!�4A+hb�'P���N�^�-:��w�á��;��_��8���=�>a�����t4���f�&��a׻�]�;/�+�뗴�K6����q��7s��\g��t��j���X%x߁��,#}�������^�[9J�J�a�2�)Ԉ)T���wV2a���gq?F�%I~pR�$� ��g�&�R�6��wp���/$�����ͤ���ߘ���6���g�	���Y��?*S)�N�}_�,�e�Y�0��Z����<�M��#,|G��;�����RF1�K-���=�$����_�5"Ÿlx��[��SPF�n�^�[!�k�5�N�a�2�&�zj��V�u 1�B���)���BGH7x|��v��0*�x/O���]�I('�z�e�n���3�e;�� ,C�/�1���.5dJ�ݖ�8�h��?�g!�f]/���:�k��;��/!���QR�Fխ*GcGf�D�z@����cu��-2�4NG��I:���"C#�� e����W"�	��vU���t��?���|�JJ�5�	�q�1#���w��p�w�Y
!\��u�S�( �mʲk���qJ�߅�,���!���e���!��ݍ�%sM��?";<D8��ZuK�	T���/#�T�l�?�/�I�F��Y�h��Q
��`0[\ܔF��M��;��N_�nC�(m�ES��3oy�dC�j�f�AT��p��C�r�6�~Nnqކ����z�0�0����w�0;�`#��h���du��"'�G��H�[�I�m�9���Ȋ�9)c�	��}���?��l�6F/2/,ۭ��T�t<�BF�ӥ�I���EN�����bw��l�Z.�7/�?;�M�,�C��a��9zu�<'z����C�y�����%�%�"O$2і�'���+iKH��b?����N;��vL����e<Kv#�h��9��*���� YƤ����V5�*Z�(�)����P���"��
�a{���&UF��!��o�I�b�p�����2���_=�����!ٍ80�ɟū9I)Փ&��`rJ]z ǣ��{������bZ�P��0jY�=������=km��c���?�:c�W��¤)��[�� �QITK�U�o��d�/�Y��vΚ�ȴ2�80�W��[p8kA�1����x��?6�;�y�0��L���ä��#.p��O<Q貣I�|�[>�KR�R+�h۞X􍿉�&Ԡ���5A�D�a՚���%��W����k洖��ݶp�}�M����&�=���#ѳDEZk_�.a}وa�Kill@Y��K����t
�dV�@���H"6.���a6|9��R:w�\�]�!�;6HР�]����J��rYOr��a��b���11?�.������E�{���W���-8O���'���q]��D��l����c%Ed�E14��]���G�����Kx�P���x@G���H��`1س����]i�֍1�2xy����3՞�5PU�J�����2_�ݳ:�[@k)�lo��u�hɤ膴.ܣ�iQ�H��ƻ
yu�����zt��f8UX/t'���2�@�j�#�cg7_�$!1W#P �-$[t7�|�f'R�~��u�}4�,׀�ta�����$l��q/�9_^����ɡF�= ^���"��SX�1h]�� p��i��=�i'PҾ��^�)E��J*ӤO� $��F�x�T�e��k�,��3�Rjx��	Y�j#�" ̅8w5BW�_�B�A0N	�.�'�n�e��L��	���{�]��1A[��B�o�l,=+W��x |��뛐���6��_堦��}�D� �&�%�O>]V�	W?�,z0�V��mB�̳oC�B˙ڗߵzCo�V��h�h+�aB��n�拉�-�(�A���c_m��9�����hieZ:�;��p��įIc���UQ4�O�L��2g�ѺFC�����d�b�nQ�Yr�5\q�����q#�[)p�A�Ŀ'J^T7~��,�ӷ�����𧿠40FK0O��
����ʀK�ՄV��a%�?�'8@�<Ɨ�$��GR��3�������umS,�܎��<��,�֘�gzl��{Վ�]���<��LM���)0�Vl�Y�<eN�����6FMPn�%˻=�m�@9\�4i@g�p`�88��
g]��x=_��� B%Xy&
tG�& ,D��x�:*�lFƾ�9%f���Z��mP�w<F��7���O+sXm]>�4��vH�!H�rT�-|�4� 9�4�+��"�GΌko!j��_x�3�|�,�u�X����3�����a�R��1�!4��ʑδ؊���dr���6�xV�i/�p�`�C�L���h�bm�̈́4�q��|�)dk[���*����U�A-Sߛc�x��?s�Pw*1�^���vOh��t܎�ѶTP�?]o��#@1~�F��C��Y�qM (r1k�ז�6�(�]��Z]HA�2.���׽<*4��?W�B����ox���\���J�=,v��[�K�*�Kw\1W���9&n��Tl���+�d��M0�IdH�όMNbM��|�p�>G*OmPpHO#��?4�v)w���8������Aҫװ���#qӞ�Mz��NP�{{G�<z��|���@�$D�3�*і�f=�.r��*3����i�^��FcU�� �(3�JՀ���g���Iߴ�CM��|����L�� O���1V����=�6�|�K�:b)ebUq �(t�hr�e�1n_CT`��/-uq�&��:i����I�nOx�s+�8{DF�;0����H/���*�(Maꅣ��e��*��l%\!p��s~֏i�l]||w��u�V,%��K459:B�6��ۂǤq���-^�n��ȟ��k�(�u"粪��4z����wm$b!T��y�'Y���C?��)�49F���8ϥ\���૓�@/�ѽ� S~I���~���P?ۯ�S�G5��b�z��h���k��W��7�;{�$'�,�N�C&�I(��p��{E��p� 2���4���CB�V�X����2��9��}��wn�&��	�ԩ��tͽ���-4����#)xR��i�cW�Һ�ځ�D\�؇c�o�l�L�m�J�\�&;�4�A�-W.T������3�q�"�%��r�9��s�������p����	G�T4��sB��_rX�Nl���,�`2L�r�o��p/� ��i�
h�B���Z̽�M��%���e�OW۹��U��t-u8d�u���~���>��5�9</#��ZiDTcE���Ƚ��D���<�xF���<���o�du{ʽ7^�O3q��8ܞ3t8�j�l�����6D���+ty.��%�>Ck�ڼ7lRTa0�=[h�W�^z��L R���2�.��W�4 �
#T�Y��(��/K��oS����Y����)qG�C� کoD�X��1Z"q$ u�r�f$��X���{\z2�HNS!��c7(j%�� 	�)Bel�#2�Ϭ�
 f1����
��x͕��`e X�O��{��g��le_60������NeK�~�e����V����x?�؁c�3N��EA/QB�6��}����g����e�A*�@t!9h��$�5���O��0WP�1a^�/���jtE ��U�W@� ]��$n�u���![��U���&��c�D[���ǡq�n��5ԛ�j@�o��Z��m�Da�F��B��Eb�g��s��Vz�k��Ď�u\�-���JD��@ � h˪�,^f�,��R����Ƚ��f���AB��.H����l�{��~-c�����)jUDG�q�sz&bi?V)�<{����!��\_*r��FfB���A�X��_ֻ��b�-7Kk��{��9�A�kW�wb�rtZi��a�<EL����4�]�(�L�_�-��xK����2G�s�ŧ��g�Re|!/;����}]2U��4P�:>`��60�u��jH�
t�EE�����\�����+"j��	�u,���z7�%KO �c�v�E�x�0ܭ��sl��o�	uE�Dk���t�[N螥䪉(�M�<��=�wfM{��%z4:�6L��v�Mϰ+��L�W'�WmOJ��2��63���h�54(]ŖZT��*�������t5_x�3��f��֔q��Q�R�e�r�+�E�vЂl\�8�����Dtk�����Bmȥ��X��|.\���,��sf ���=ڭ�n�~&���\^+�U����$�O��c���ך	�mG���l\���9A7�uuF�mo�B;f��,���T�A��{W���"qey)>����^ie�j��}*J�,����=⼴�p��5��(q�g��%��*a\��a��<��[e��iӚf==d�`C��8Ҹ�Z�	��e�ϙ渝�q��ޚ7u��/,�%��l�&�D!� >���t;���9���� ������,*����Ѡj!H���;p�lofV�=�M8�(�f%h9D�xm�O��{U[K��lFnS�Y�1�!C[R�H��+�l#���ȧf::4ȸn�m�t ��v$���LZ+�!�r����4�]�q�z�5g�ڡ2<�@}I�<ʰȃ���������!S��5�|&~�ႏ�sX�(�.��.�"�̛f�S�D��,2U���;��Y�����ȥ�@��Z�. (Q톎JW �=�
��>�O7n�7����T��R�����z���8Y����k���D4@VN�T������s�G���Q�&6�b�}���i�S�n1MH,����Z�"5P�eX��;%�I����A�ĕ�i��PCȉ��$�Q����0 y9�Y\P��+�Gn�I����]	k^W�����Qݩ�׎}#N��E�)��t?�o*�Y��_�UP"%�^����E��"%v�$V�a��t���w�Z���x[SBD[����I\�uR�}9��?�<�@m��%c?��]*ұ�������~�z�OMݣl�+�(v���vNT��<�F��T �3 L�J��)ΡF<d��v�Hwi"��IP�k�]�Լ�M�����c��y'�~��dV���	�/^9@�5*����3˧h꿫*�����#e俽;�q�P�V�����R^Ne�Z�üo.4!� y\tL���  L�̟�)grT[L͐a����0Z�������=�|Pty3?���|c=�Hh��y�ҙ�P�,��w�^��L�����Y��$8�ΰ#)�ukT�ÿ�=��$�I�@( �35:�n�S"C��;B�av� ZE��I S&[.��m`	�	�/���O.!��J��M�<	�3�²;���)V�ΓI����H$f���"{%�gs����%A����P.�sr �#p]�݈�7�G*H�@wc�J<54E(����ֳ҅�\��2}�l�|�6��3
dP���z�{��O��-?2*!����	�
[�W�'T���hw`-�3U�� R�]��a�2D:	�Y�ና�mLm��L�z1^�y�uv�"�;���c#-�����U�@�ӝa�^�S�R@/,�&
<��M������ۂ��x�b�����_�}�͊�:>�XB����5R�"�a\{�B>�������rMV2��/��%�X0�'w;�9��Ump�F5ó�u�����N�03�)����蘨0d:�;wSBZ�:���O[�fg�����b�$�A�n譕�ٳƔ��)����"�@-��4tlc*U/'�&���K0^��������0�7ñ�R�.�Q��lL�%��T��M�~�S��Z��s&Y+L�f�9K�e��_|Qz��K����+D�Oe~h�nnƖ@ULt���4������9�W!;͠O��$P�v�z�꣙��6 "={��\�ѕ��w�e���D5ڑ�`�MT��X]�'q���Ĝ;	�k���nkE)}��f㌛.G�6l����+mqm�=���SY�$��i�	z��� 2Ov�I����8V�#Cݓ'SWv��� {�-
�V�#�zq��A��V����^��_�=��r����
����� �4 ���<�$z�4�z�W1z
�̱�
�0�ϸ��.��$(�:�����+�"�ji
��{����y���:l�c�n*��K�3v�xe@Eǟ��Yq�eE�{��_�WT\v 򧥟ޚŸ%1n}��8����Czr�~���vy�[8��%8�Ǳ��p�yhǍb�_,$���J2��}�����=qQ1h��0�r�����$3V����`oP�L6��e��4���LS��z��R��A/w�++�9�s�ÇjY�+��S��^ߛz���u_����X�h�o��]���]�Y�'�r����K}y,�X��G\9Y?h����0�P#&C�ƦM�@��Ҝo=
���P��F)�Jwf�~��BU����h֗�|�>��~�ȁn����m�7�v�����'g�R�Q�C}82�ۄ���-U����Y��Į'6`&	�u�a9�$#��ͳP��p�����k'S�M��7+^�t��)�u���=�Sm�\/\���Y;vÛG��8cK3�b��:CΥ+]��0���
����bi�OBZ�� �ڇ^��[�;��ػ��D�o9����jL��B=ߏ�t������\����&�����_�K
"�u�����?Y8L�Xʚ=�am�H�L+N����C:���U�r��F43jO���j��!^����N\݉s�JT��+�ƒL���Wᦜ�L(�����Op���p�:VXT;�G�C�֙���کъ��*���MU۹�#m�y�$�c�)�{�B���}���IZG�\Q�<�1��p���9��Kq�ъ47).mHԃ4�j�t0�H+-��D�`,������E��X��2:�q���S0�{}wW�'��~�F�b��[�b�������N��1pT	4̸�f�LӢh�i���[_��X]�����,.��2d��3�@/E�E�`�&�)@�8��1�S�$�@n�ƶw��2�8P͈���ς�X(��jz#u[�@R�pd!KA�b��݀E�
��͙F�Ԙ��T�� �����d����ʢ�`�h̍�.n��ݧ+���#>��bL��Zg57�džM=y_&�.��	�漏�V���~� ��t���<cN�Mpjj��Za���<;����;<֕Kی�فUV_�N�1( QI�j�ҹ�=�:ط7�}��;8�O�mCB�I<��
u��\Z��ԛNv�uj������!d��	KKM�<�ήY�nBt�Ty�c��v� =o<�C�R�����gbB��&��4]uQ�Z�HW^�+���4/���U'���F��ht
߈x�`������������rE���N�51�(!��}� \h���H	��@�i���T	dT����M�����U�4Qv&��v_�����J���s��!n�j/�Ƴ&�ڝ����B/`��!n�j;��Ѓ�+�_J.����*�G�[KY��6�6!Qc:���Q���=��Tv2@�F�/�X�