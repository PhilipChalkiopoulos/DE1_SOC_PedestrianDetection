��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b�����:��@��K����[j#��������њC�2��}���Sُ�7l�l׳�.�SF��
���qmjlH�(/���ဈ�/ݴQ�r�1���λ�_]Q�K�T}8s38Ğ]}AB����������/e�~.��`�����ĺ�w�/�UT�z���a:�)�W���_����>���P z:d�Q��h�
��D�!���n4�h�Ao���iH�zv�B��r�z&n����.Sf���SV�a{Gp)��50U�{Lg�FQ��z2��x{�>���_��%٩��å�d$w9\oɓa��"@{��X�Eല8��-����ȩ�J ���g;��)[��d�����ߛ�Da
e��#���4-��[�y	�����k�y������'	u�ͺ>gz��DxY���Ϫ�67�jnʄ7����W����9���/��Y9��/>��N�u���^z<�M����z���O�,X�0��5�7Ֆ�;./9��T[w�R@�m�P�=��lL�D7^�#^�e���������µ�Q�#��E[jx�♤&�d:��@f�?y�"����d�QcaFK�t�V�)qb�d�ze�x��$��|�� {�9��m��U��j�x���7���tM�C��9'�S%Nw׫�'?<��g.o��k#� 3�i^�� וӰ�k!N%�_���%�<[�%xoQ?��A�#<�_%v�w@�6� p�Ty��  �/����~T��U�}�Q��1O�F��k��7�U����lF��ɛ:!�\	W�z/ɗ�G�me��G�C���F섰��h��y�J8f�K��+�-��`���v����HE�
1����
�l�:�ǳ���% j�}RU��L�7^��x�(�y&G�����?˞S!��K-�C~��﷡O`uq�Zу�LG��W����MMgp�'���U�vSޫ�%,A���p��ui+$Tō>�.�}���������D���Z&
IN*�4:��L/�Ԯ o�[��ɵɸ뫤'�w%���6l!G�nɆ͏��&78	Q��A��S��m%σ�?�]J�$���#tUG�̭
krG�-jPp����j�����°�J�,&2F	1w/����OƸq"H�q.��pt�g8ٮ�9����8W$�p�g�$f6�O�8g>�ɽyL�L�$��6��7.FS��'B�3.k���_\�3�4b���	r�/��P�� l�hZ�hB̤m���s�:T�&����H��~,�AHG0�S	����Y����?9J,6�5 )۸S)�.���,��uO�T�l�u�^�?7C��{�������!0�G�#z���Ee��k�t�e��{���&Ј��q]} �h�S��Z��.v�&���g�W縑rЀ�k�A�w���!�K���*��Ո2z��^j��eW�EM��g������j�ID>6������E�ҿW����˛E_��L��2x�QXBO�� ��E2�s��Uw<��P�w;�
�_�8�e	�ˠ���'d�b�ƻ,w[/x[�5%5�xr>-���>�&C��Q\����y7��!C>l��&��ϯ�R�Hg�9�7~���yj����HF.|=���x��p���k���5}��,����s}����U�V:�Y�ta�2����?��oK�q���,ou�$���`"�%�9FsO5*�>��齧L���>�Da������¿����\m�s�
���!���u�ذ?�B��*���� c+~Ĝ���쁌���}�]�`�2��#u<c�?�R����������H�+��Kq��R��)�P iUEX��{Φ�a�S�	|��{(>�fO΁K{�L���*�ѫ�5�	�Xu}�.k�@�v�HJ��e}�Wy�3��]_�o^��Us�~�~G�<B�j_#�اr�8oSWՈ�"�`I#�D�c�aQ2�r�,���X���$1�B�M�!b��w�ql f*S$�Q#�r�۰cj~��H�<�����o��쁈J�C"�GS�v�Qu�ǹ�!�>O^�~m�����t}1�8��&	~�\����%��8���Dm�L)h� (#��B�tA+���&��Ȇ�	�Pz'�(�9v��"������:Nea���q��˫��j\*%W���5g!|�? y��bc�qNRi����2C	Y�=���f��^^.�m�0�ݥv������?s�u([6�˸}͛�F:�؄4r��^�&��I�L��(�2}2��F�kO���]<F�_c��}�̈́�87G��7�r=��yNF[CC�/�J����W|��