��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���jl�7�x�֫����_��aoY��?#��#�r�m�"R^F�(hb=��pt$��e[5�v� ��n{L�x����o�x�+@wM�ca冐堏����D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�KW�UHսQ�����_>����ȡ���ē���a飏5���� ��9o�\y�����{�q��"�t��;�$D���e��>%X��:ot�k�k
vk��S����A����9��}w�9��"��ȳ(Ym�{^b��|#��0������Rah�֎�Z�� ��7�:�o[KquA 0תO���К�:����˜i\�|�����iBn�6Y3:�ȣ��xA��=*�a�;59�M�&e�Բ�p3D����1�]��-�i�)���m����m2���0���bFO�����hX��6�#���t�7�慥��MG����m���(YA���O��kO��\闖:����5��mT�
5��V��y�iv�K'���<J �w���Y|;�k�N��,�������#��e:V^족�j��r��&ט|�;����L,�X��N� cƖͪ���dB=yk�O,5sT�b��If�K}=L���Q���0N��嘞���ЇuS�;�5*s�>=oW)���$�YzPsM�,y/��R0��$R'4��P�pEo�gat������6i�z���|�`;yJ��%�^>w���:�v9�|���D.�F��&D�L";=�L����Z�j�$����!je�*���2�b�><�+$!E�e;["f�	:��^�e�_������砅�v`�[Z���-�=vP<&��oưG6�k���`o�W~հM]��σ�u'���N�ȑ�?�ۅ����s�r|����7�
0�p�O_�6���$p��>Ό<��M�C_����>�٬��������@S�v�f=Q��1�l�����$Z*��<��[��b*F�ɒYX����ſ����B5��Я?�K),}&k���B|�!5��{n�c������6�г��<W�Ģ�Lgw�W��,��]*e��s���Ճ�'U�%}��ً����x�w)&7��.��̎�F0Нr�l9����B=j�:}���A�%]�'��9>�{� �������u�L(�r�ND��&F�p��}���;�p)c��([Ҋ��vm olj#��#H���{����#��;�)"�r\	?Y@���փ"��bJ*?�w���t����=b�>���V��
�82�5FSVŲ��\��O��{��1ݤ5��7#j��%�T>��Zy�U�b>����3k��/L�ȉ���erJnL�3�FQ�����&2�"�7�hWa!6��Q�f��/P�dc��x��[�m{���"��o.�3G-N6��f�>�BNC�����H��Gy��o`�H^�3�EO�mɒُ��Ւ� t���:��&/*��
�*K��q�<�~O�t���z���u\��+%��E���j>�D�������������E�M�tG��kj�~@�g�%_̅����-����+��q�޺:5cP��Ck��@~����������	�.�T�`F��C�	�Q%������fQԅ 6�O�X~�������l;u��]>b�G���Ë��^Mq��$p�[�c^^������m����u���FB;_��96��O�*^�'�^�{$��r<C��%��I,ƀ;t<���ӯ������m�i�Υ�{���-��1�% ]�[�Semf'�4C�l; ��HG�p&L4��9�ZrCƏ�
ɲo'������ڐ(�Bu�0�E̒�B������/5���ߐ�����u�Cy��"yg)�ߏ�+ �&��X$��7�ŀ��S%�>��C�����������a��7ـ����LJʹ���RI��{kp;![8'$��SԳ��?��?ZF�=��]�K�2m�؜��!����'pH����bP�A�5�Y����۝4yS'c�^�;o������U<		��D�s�]Gg��(��r�^�ox�^��}a��������s@`�фCw��5޲��|�!���$̳3y�=r�������Y�AEͨ��3Di�7h�}�5���C,=w3<oؗ��� �)w���AFIf�!	�L2�%/9^؍���$��6�J~V3(��LZ^�$LԮ�ڐ�b�U�\&��Y����`o��.�N�[��ϛ+��+�sMSɈny�=z�K��%�[K�`�	7����f�q�
���ӝ����>��,0-�D��w�+m�������|�D�_�^����r~_<�Vnr�pQEW�B'jx�9��s�3���.Ͱ]6�u����Y��s��K���m��Vjo�4q�W5c�c�$T��5�/�FA$\�d��H�R��'6�%� J*��&Q^qe߂�9�N�y[�~�Cw���v�_ۭ<A@X?	��c�ع�p��|��)!�3Vc!+ S�)�v�)��G$��l����:�+i]�}��V���waby�<�j%��/F�,�d�O����S��J9�ƚu��@?#���T����A��J�b,�8_�d7-�^l���� �Zp5���
i���F_�'F�0�8Ѝtv�G�-VxG�j����t\�&�U��`��Y~�<3\�AAfw�^�>���j�wT�b�_��Ia���� u2{�?�$\�M~3ǥe��p"�j4%4 �_`B�N�0�Djb��l��K��)��-bs�e�� �[�tfc�rVM�>�ĨZQt�͎���A�r�	ч`�|��M���+PȈЃ�����z���{J��B$/���2FΡ���2��-/m��w �}�3��]�h�h1Ȫ+Y����v�<���z0]*ܗ�^	ٌS9T��Me�^yLue)�>i����͍�F�c咳�p�=�0�����ݟC�t�Eo�F��q?�^�n���w6>_�)�&A�<��* o�y8�y���E�P��bF�X�r�����Y��-!�=�.L�86L��ܼgV�5S�
',�?p��M���G�T̗Y�4�� ��)�xi,Չ�Ӻ|z�k�t�X=����`�3z�8F	��%��z���Ƶ�Iso��\l�+�?���'�=^7:�ߑ��?CoB��-}�Id���xIq������o��@2��6XEjaz��q8z��d|�U���]k^F�J�K�M�,��+��NZ��B���� 5ֆW��	����%|䤺�����+�s)�!�H��n`��1��4;#TQ�vѾrDF8呷��[?޻���JNlݣ�Ǒ����s�}�O�|/��Þ^*t�dN��Lf�T�����J�����8U8�)nR�\�i�'�֝h�m�r�[�޼+{�)��ޑ�pSƈ�`ç�y4�D�am��lt
��M�� �9H��u�+QlD��	�&����*�����q�k:c{��<=4Bscp�E������YG���<W�p��w�Oj�x�E�*�G]dT������c�l�ׄ���:|�5��	�BaĎCd�C:�y�(ey����ε�4�z0���!�WC�).���O���X*����)6\�����	��a�D�+���5R��'�j�B��`�˗A�Dh�e�` ��]�mT�_˃!�r��϶>�\P4 �
p�7�U,5�QEQ���En�	{�=��O�����lt�@r�T=�͛޻�ȴG��&.(C~��$9m�1�}��R$�	Lc�+0�����r������	�x����R6�&���b�Y��K���F�jy����r1�C�M��ٔ/ob'}����U�D�4���5ݒ�7��L�t��X�CO��M�-��<H���T#u-��L��I��/��s�J����)l�����$�q)�1<5	zgA�X��!��ٛ�|���Ѹ���m��S2��b���;j�o��6M�`e*Z��(B���:�s8�58)e�]�uM�/���DS�g��5��$a���������K<
I��	��:Ӏ��s��x��ZK��ߙځE�Ϲ�����`�S~K�'�����=��m,wi�G�b��I����Q��=��X�3�F
C��0\��d�\A>�e�8�I�!��+��MU�
�q�,&5K���Ss>�V*N�f�ʚ�x�=�i+��bd�3���dB�A�X��'֣��[� �c�@�ג�8N��ĈY�-��A)��m����	ɁB�E���[�ݯzk���F�
*-a�V��f�bk ��0�dU�ݐLVM覑}�G��M?��8�pB���Q;�@ӝD_qWx�4H����S����A�f��s�p��.}����Š�+� �nů,ַ�J�6�<<jVo3�wh�����m��%��a+V�_�����`�|;�4Cm���
�O˥���?�Ç",aj�>�7w~hצHP���>)�i �!�@�A(�Ģxi�X�c0���Ӑ*L����� �>��^���X��UZ
������(������jr-}��� g}��X'��b��N�"/}Y�IB�zn*�ޫi9����-���vZ�b;#m2�`kr{��H�OE���y͔�� ���p�\\�ɓ�4{Z��VKO:$Y	�F������'�h����5�:H4�`9{l�R'|k���ّ�3�>��J͊9�7۟�|�Wmm�f�'!7�>l;�J����0͠{�b�R+�"����-��6t�����&)�R���� .�*�I��LB�]d��$6|�
���hn��⁂i����dL�	�`{�Ϫ`?�?���B_����PK5dBA��D5�?괍c�Y)r���3u��`	7S�$�o��_/�W��_�dޞoÑN'gQ�����x�Ӏщ�,���N���;�#AKSX.���k|��>3o}J��W����Y6�6mm���`/���w�Y�0��&��pO��[�,$�����C��T{�P$(O,�K�H'|�+:����0n��03a�T����\���l3R�����%����ށ��Ⱦ�(FQ�+eP�ܰ;��@|�R�gH�E�c�P*E��*��V�QE`ܦN�M��Ӗ�<S P�cS���dҥ7X/Y<P�ۗ�DO>��U�}
�v?�h���}��=���"K���`�Mk�Y �Ƕҫ�~X�8t��J�t�d��!+��Iav>��j�ct9bT�ߚ��d�y3율{RT���ɵ�rb b��*���ri{�U�Ǹ"/4��&�5��!�I��Â����/l���[��*����j�`��Xhi�����M��s��֘Y�5�+�sL���V�S��h��)����͖C��{co@�-��X,C��E2���Z11w�Z;Y"hW������↙�u�(c��qzL�$@��
>�#��e6$QMQ�Z�
�ִ@X1�]b�}��b̦�1����mG��P�P���,�7�<�z2��ȉ�m��>s7-��QG�w���?1ӽS��"�����ς	�*�}�k�H���7��ClW����h5�&��S�[�{�`��"��2�������.��ƌ���?��%��K���5]A�;=r-6#��c�,zo�mM�h���ج*�S%Ͽ�!gl�K´$빢��W�'^myVz����5�>��qa(�킍�������"��I��K��QLb��k�A|���?��t��y���Ų��S��z���J��耏�v>�|��[���Aq�X����b�� �ǲ��[D�(x5��8�a3����M���	ϝ��3Y���
��K�,�c�nQa���&�Jz%�-@5��%����OfI�r�����j�	�;�\�^����2�p�T�J�[�@OS��{��E��ƧTV��(��!���H�GjF!�8��S�;��te��;c��P�$���.�"8,hG\�����*A��	0~,[�\�\gW�:X�yeF4\>����!��2��0��V���fs�-@���u�-�z@���9R�K���͑�� �X�q���[����c����s��Ç�d}�����g7;\r�x�����WѾ|CKu˶�������?��oeg�h��Ϧ=�`�K���P�����j,]i�9d���4��Rm��&�aS#ª�.���~��Vj@�6: �_c>3�,ۧEtjK�
I�K7_�1׵j��c�;��F5�[QJ-���ڰ͎��!�=$�5 -͚�tYߡ��.XK� >cʐ�/�L��������h��j��Pn��(�f�X���4n����@�o� ?�i�kW�ވɅt@Γ��%�w��zt�A	�h���99n#�K��ޕ	w}�~_���4�L�)�xj�ڀ(�
��Ԫ3��鞗[�~�W����Nw{m�,D1w�'w��'���B�87	���̹|�!��R��N�ap12w_Q\U����QǆP
�*Zj�x�?G�����M�{�~�G�
r�%9�{�74R�]��	�u��o�g[�0"������ ��Jt�Q!�)�?�S��܎��Y ܈�p�h�6D��w;�lG�%�l*w�K&���-i�0]����J	p����|�ʙqt�,(x��[ق��>\i� �x�}1�Lҧ���M;y'y5:˧Ię�mq�zp�����o"[?���N�����J��k[�3��b��C����b��C]�8.�&���j�j)I���U` �0��9��aB�\"���J���@Kv95�ڈ�������/��Tm���7�Ex_�"��s0Wjo��D����
"�-������
�*�sf�j����Hd�^D749қ��s�����,I6�ͬ����b!hќ15���[���q0�ua ��:8�6��N^`^��J�`����T�݉��y�����8y��<6������q��
T���J�̌����ZeL����6ɚ�~�*���>�P@ǝ.o 
U]�g$k��[�:���a�֕�ew
Ku-�
=�w���ӝ	d�P��z2L\��a�,�_{��9������7s��Y,}�S;���ԋ��!t��r��ɚq���O
��u����S t�NH��""$f�&
f��p8G���x3��w��t����M}&�Ib�&�x�H�]0�A�6���\�*����-K5j�Gb �z�x~>�U���j��Y���_�WCfk}��`w��������{E�?h����|���@�2�u��x�XnN�����q�3\\ëT����es@����;thzߎ�@�g��y�s���oP(��G�9�4M�?� w�`�I���UKpC�LP�&W���*B~{ 7���0	|��4ſ��A��]}>��[�_t�
���Dz �%���v�\�����R5�u�t^������ql	���>A�RI2�%�N���@�������ŉ�&��0���*`Y��:$�3��S���2w���l�j�,{}��6���H�u\QE`5��D�VD[m�S��:p������Y	���1�1\>�k�^�l�|��t���A��KȬy=��^B�d�>�Bg�˷�P3J�6���SJFx<Ԏ��c�g�O*B'{4`��[�b���A�Ѓ�=��B�����ҵѷ���ΛM}�>�������JKORK�M����g�.��4�\,��l�:�O�e�<�P�$\�h��#ݠ�h��QMs
���P������:���+L��c�M���<�1����8&��I$�#ޞ�j�������a���"2��P�lhT����FҬ��R�/��B������� �$�+�CƱ^w\(&�1쿴%볡��e�K�ե:�ACe�l����*���˜Z�n[2��@7�+
�1�{�W��:Ұ>��򀥳��#����"#z�YO_�XV
:�f>�(��q�Yϵ��n_YvÿJ���r	zW��Z����Vi�6;�ª��5 �hy�z̩6�]9��N���.t4�,B���}��BDz�a`:�Q�� �6!^G�srp|-�`�N�ۼ-��U���_��G��!�?@�Z��Ӳ����da�˘�a^fS�;җ�E�a2Q`;�#�7\��Y�x�R��BL��O�ճW�U���1*u���Y�%��$Qx:d�ݤ!�Ł��BlF��p�f&�d ��K��Yki=�E%<(��(Ɩ�� �C�]�+;�;7�S�8mԑG�^��=��%�3A�&H�a�f�ʺ�.U��ш��		��Z��:ch]@rX�vr"�mPA�S=V�I�(�t��a�c.�i�A���è�"v	*��/��$q��ml+C�,��Z��~k.�.aO-4h}gz,ӫ�R�Ԋ~qF~�������oU5KK<��5�����ف"�
H�`&����=�n���o�9����BJ{Q�՟��/ ��AO��g�^ ,�D�z���}�'�##[/zW|��,W��3�G��U9�Q�V܊,�䍉UoLY]^�d��T�>LOiM�(]��?�5p�I�n}�f�|��T�	����]*���&���9��Ъ�u�J\W�b�Է�ǭ��Ҵ wW>:���t)�&��E���>�"�_��1@��-�z�4*��ݜ&��W�7p3!�ź�h�#A�*�*�c8Į�������g�Lw��m!X�b���������M���jU��$\�cK��C�չ-�G�7�Y��dݶL<�Z�4m<�y�~���K��)y���UC����<ΒD��b?0�+Kd͏��zC&�p3OtW�� ��V�:_�jćWl���o�G�"�e:��/�����������[��v�,4�ǐ#�%������g�`zZ�0��	�9!���x�9S���۲����}v�(5���躮��曹���[�[��bRJ�e�2�'��Eb�Q�n������l����|�R�����kL)� �M�d�k�l>ߗ�1 �Ͷ� ���ك"��s�ї��s��p�\k�~x);�2���W7־'�B~�dMX+ƶ<3�( �߭WI�7�%v��YC���Z��i��ت!����h�adb+:tj>�/�"Ǳ/zj6#����Y��c�q�8����(��AE�E��"����s|�SI��o��P�n���ގv�Ų�H/o�A1�~���k�USI7��nd̢ם��t�(�K���n�!1*0�ȋ��:>��b�A�� �MA�a /7�n'��,��Y���<���@URi����) ��y$�[�<���)E�"�B�����^��|$��`���=pWK��kH����2��D���>�Ȭ$$\�q�W)c᪲�",�G����`}
d���wqA��m6j_�3���-���7j`�	c=�2�Y[�my<x�)n� l�U����w���1�8�cI�L4���W	���X���8��L��[��6ϠÎ�ˌ�����F&9h�}�q9V���z���r�a�r��c��Qo�9,>g���-��|i�����t�����z�$A�w�����QHoU-V��Nц`Đ�0��� �ژrTM�����N0��3*1և���"��*�b�)��EE�3T��&O�s�XU~���R�T3���w���aΡ��]��!������6~��'�18��)8�(��n�F�QRk\��&�3�j��|�h^E M'�ʟ��S�J�o��7��ۑ�e�ƍ39�~a9�-M엦�H� ���c_ϋ�>}k��:k}������2�c�@�ME�p�N��}�Å����Z�FG�~�ά���R��$~�k�K�-1�r^�668�'��乭Ci�
�z8xM��+�)�	�W#,u�Z6{��tO�6�a����@�7d�c9:?9�p\(v^�"��s?�x�	b��gi^�VZ��KkN��=�K9��R��x����VI��}sȚX�Y�,�I��Ŕ��&�����j� �~d ��G�*���(:��Y�.���céR�i�NcJ�5��`���^7��mtA
��)wZ��"LfE{/�B�l�nٖa�v�G�'�*3���9Nt�K�V �V�]O-���z8������)��0s�Y:@��m`ߤ�7�A������QθI���:��VN�G7c��F%Ѧh���O[a ���_?��	���I�$��F�C+�{���IMq1F���=�5��ϐ���]�)�/�C|��XѾ��l%�j����}�m�c�{#���.��ZGW��!��f�#�Z? )B7�x ��r�?S{ˇ�3J���9���	���!�&�|��싪�-�G�3\Fn����)`�B{��10�s�d�������'R��3�S9��?��Y���qUs��ʉ\�_6�S�i�׿�i0�8�=�S�)�+���ʌ�I|��Gm�9�	���mX���s��xb��A��7�Ϳ\�ln��G�1p#��R��H_厳�P�4�&L�+u�
#���:��ρѰ�h�_�<�� n�R���-�����c�`7<�7���s$��vF���e�M��3�P�I�n��.Z�Fsi����s�[���M��5I��E���.>�T�5S�:�q@�*C����Jћ��+����GN%�Q�!��?���|%#=bi�Cd�2y&�P���+��)%l�`�K� ��τ¯��avfȅ�!��ިs	A��3�����gRj��*j�H�-E.8� �?��4�`����r�mF�M}0����[.�� ��A���18��w��)�����������1(ѵ���d�2��-i��"���Y�~�-������(�+���"]�?���`��i��9��B�n�����s���%�̀��ȟ���I!!!�z]�]!2�{�(��H�yDG�I��$j���o���M��8��!�����a�7���:�AY�@�߻���N����ZKa��٥6�b�!A��H�@{Ѧ�!h�͢�-��{�!.i���8��R{���L�o��-g�74�����vk]���[}cNz�dB�AH�y�v"AP���7�*�o���1�~�j�|۵���Xqk�����g���0��MB��O�ȕE%/�I��g(��10F���.v"=t�h�J."��J��Kf�O{��=s��?�X���Z�d�'|78�94	n����#��1/>�]�lހ|�em[G���5Tu��[0,Y�r�Ϡl"L��������F��X�!�(�^��܌g�,�W�p|��Ѩw��Z�c46A/��P�Z-�(ʲNcy��Шg��^NCڥ�E��|��m����x^���|־��Ys:C�h�l��qFɽ��u)Y,at�(-��)���J<��[��,�a����vU�6���2J�68CkB�Hwc��X�ܚ�3�p5dq�`��\rz���?�SZa�[��ܤ M��=~����g\��'p9�{-��z{�m~��紼"N��w��p��Ȓ_=븢��ݫvφU�5��MķS)�lμWN;e��������X�c�L�tJ�S2tZH�Cw4�3Bͬ��`�zB�cQ�_���[aQt�l��v�⭀�q�Hপ�%^�����w��+��R����A ��j�q�	��ƫ�i��.ߕ*ݣut���ip��Cէw�ő��z��l�};�*�6�jj�g�*� �Ts-��M\�B��I�Emw~Y�}o�%�:f���zM:��Pkምa��X���tM��Y�1zq-Bk|�DB�����j���8����j�b����5��K5�K������]�hmT�LtsOu���x��x��Z���#�!���d��#i�)���]#�K�R�T*p���&Y��Uy�\Ń���Ro��C��K��l5��(���_�"ve��/��Q�+�g�����ԥ��?t�[E�)�R�
�L�L�^��]�q3�uXW��I��y����Z��f�l�xSa��h��#.�5�����#w�ЭhDl����[�kY��Պ�2L۩�.�H �Z~��V$K�����̸{wb�t9$ȡ
V��7�� |�)M2o�uu�ٳ�Me"mrzi�6�O(L�k���ʕ�むp.o���.����
��������w3~ܸ��"�R���-Vb���냟 ��rײ���J7�@�� �}�M7��>�I�P�{P�`FM^�,��#�[��뛣�@?o<8�W������t!�̞���a}����U5�:W�8��9�߼�/��Cn��29te�-�TX�P IV^�J�c[D��. <eQ��g7���JFʀe�a-ʢ�P�}����μ�[wn��dֶ; �;̲�m�:�+���l����*B�oU&,�'�$\�Q�HXc��0�W^����)���5<�hR_8#� �|��ѥ���+8m��}r�噗i����:gx-�7�R�Tl�q:ǯZ�S:,��B!�1N�H]ϧ_ ����R������?����}��gy���N1���Q��BjQ�U�p����Yꔊ-��C]��+҄ti�+I��w6"�߄�ᗌG=�^��2�ϖݔ_A,ٚ��+
8�u�^(���:݇���%���]=RUh�f#�N	é@���41��T�Y�����3��9��1����B���mB�p�1��nS?�P��s����M�T�[/&�ECި�X&ܮ�@�D�VY����A8j������&�'�2_=h[F򶌼46~��c��O�B���*1�+���Fg�� ����t��, u��i��	�� ��Oq��!jl�B�������c�}�k���ǌ<�S�o��k��1fԑ���P�L^"�-�q��K�􈯰����݁z�h��e�s��" ��	 �ˤ���IG\�-L#�v@5��(QLQ���w����i�0^s20���ג�Ig���Pw�uk�V��!��ݾ8 H�ޢ2{I��A�!�����������5�[bXY �w�Cva���i��/>_��9�"���J:����Gp��_������V��
��R�����O�����DBϜ�_�����dW��ֶ~�]r��2g��b�5h��ɳv�,���r_y(��y��8�Wt�)�� gw����9CZ��BY��	��D��W�AQ�&~-�_+��wP��M$�ل��3�<�:�y����Cܟ^٤��BApT6o�CMR���9��C�~��}5:�mn���9I]\�(8��)HB�-�j�K��Y��z��x�v;��͌.��!����д����B�k�`XGP���1��ƴ�5aD{ ��8 #����X4���:���^���x��L�q�F0J������#т�>Ք�%��+� ޟ��\�cB- ���쮞ژ:{�L����出 H֋Q�e�=�15&�tJZ��h|t�(�u��H��0�	�x=��sL�L����3���:�e�h,�3D�𼂓�
|�>A�y���	O�JS!P_�ĝ�J���\���D.,���u ��S� ��q��j����x�L?m�Z*�_v���}B!���c��/�ǦK�M]��n| �Gk_Jw4�hح���K�n�x�y�T]ݺ��.�@5#�<�&
�n5�",�58�u�8,ߦ(t�Y��h����x`�piV;���EWR(,V�Uqȃe@��R`^?I�Փ�el�(1T�F�Avߔ�����Y�m2���Q�c��m޽M�#=s 
`�D�@Ao�}�ߕ��<�;O��6��w��&J7�ɑ�3�#����s�`�(�C�r�� !�F|�4|�Jݓ(�F~�.V+��+és������`��A�M�ǉT H8���]yϚ���i�:2�-\KJ�l�s7��)��}����9�f�h"{$ _�&�7/Z�o�y��~����O
��3C�n�2ۜ_��[崊;]�/����,�QUY�ݰ�Ji��v�� �j�39;���\�V��I��-�i���ux0Y��3�?"�� O�/d{sڍ�%x� �;�ٟ�]VK��M��v�/����a0T3-��}�$���ġ���ߜ�S�tT��V0���e���ZF�%���[>g����x�br�|���l.�5�Fs'Qꁵ^�Uv���Ǧ-J?b~�:-^���eZ�;�[�<k��)�����t,:�P��p�B���z��%��3�'=��I�n��}��1�d�`E�%u�C�<jE��bA�
� ����)��i�΋P�]�l�)�w"��i[� ��ȼm$dH�^|�U5�^�$����8p홋�K#�ן�lc�M�����1��J����R��������^��	r|�c���J����i1��wO��#ח�X�����E��i�	8�
ﯥ�?�dB��[�(B�����_z8Jap�_=�����2)یh%!�K��k���!��ъ4c��x� ��v	�/l-�~���,ld����sz���Ʒ���3|{qY�=�s�1������P�Rm�!�ٯ�B���{����V=�2�Cƪk12�����/l,Gf�e�:t��:n�"�կ�sg�u��}%��课O<yW/:����k2�R٧��m!I��a�\*<{�&��=?����4�L�
��p�.�CIly�ZA���ߕd�pH����5]p
��n�	'��-GQ�,�&Ţsǻ��5gD���kJ+�j�.�cvsms��>f���g�p�!mU�+�hۖ�$��P�Y���bI\oF"k�Ǽ	��G�Q��`��;��:a�[L�8zHn^=����H�U�6�-���ZÝTZ/��X�E�s����ھ��T��������	���u�M��Q~&����2d,�!x	��n��ˊδ���q�4;���{h����s剾�`U
��=2��L����G��J�1��-�{��9��2�9Qĕ0���r�V&�Ѵ���v-�ʩp���0�~�_ �Ƿ��Q��8��:Ԝ��Qv3����S[��_[6���T�<c� �������l��4gRg姬_���ΗNȧP8�@1Jx�"�ɡ��h�;��򖥘c�1�ۺ�n�1b�V��m랢q-j·/�,��E)��bGl^g�|��f�"b��>�-�N��^tB�I�����\ky���J���"$Ί�t	z�t��G��	�&�E�9�~^ QH^]�T����_*��w2��IR�ԲO���1�br�����Q�W8`p�A��ԑ�=���U�ŭ�L-	�s>����{����(�P�1��C�eȹ�˱X~Ѹ�ʓ����.�o�fv�6�?|2ѯw��+�9rƶt���}]G���q���rf�4��.^`�f� ��c=��Z�?�^�YF?��S�E[j4C�������0����Go��i��n�̵S���煝�B��$m����d!��b޿z57�@e�H>R*ūm�$�Y��'E�S#�0䜋��e
��F,E\I��/O��꾈>�����RDɹ��%05@�{��_K���^Ӭ���;��/�I07��|/�4
f�=f^�@�}����� dA-�ɉ���LeH

����>���\[��Ĝ#�����8̀)̝�8�GY�؆���[1M:Wj�!o�c%Y
���)xKt8�V�vZR��Y"�]Q{9unN��9��_8)���x{_�qEA������Ҷh��/� �Nㇲ��&˘��c!��-zF��BMS�9���NU��l��1��6<����y��o�j��x�%�}�*N���v"_��
6�p���]��h�Q<Љ�ڡ��V�=���yz+���ZW$�$�^+zN��j���i\�]��Cb���$zZ�3�I�ޮ���S���:�v�2T��j u�/>�`|M���וG<*��-`XE(�n}��YJ! pa|�9�r����Ût�e}.)΍����x�-l��׫)KP��3������daNY��CJ�!�b�o��Z��It����k�y��/Π(�K��3�O[��N+B��^O��[����
G�!q7�	����L\ȡk����S6�lMr������UakXA� hAw�ѽu���3U����g�rchW��~<.U�AZ!�y��z�k}�M��]� �Ă�U&��#σ)r��B�,�s�n�p����=��o�W��njf�N����)/%���)�?d���1�����l�zvŲ�.Ĵ{��π�p-#��C�%m�Nj����>����Z��q�W����}�J�8 �P���w���^��om���ԅ�ց6#��T�6z���A�(i�}qLW�G���I{z�F���Ώ�U�VK׬GI�~'�)��.39a��K�Ԯh:�- ������3(H2MO
l��	�0��D���Qq��J���%�c:��n�|;.C�"��rأ���P}xJʪ���hF��ZX��'֊�L��3�!��%9������fk�*����5�2(F3cC��bݠ/��r�WM^;݋��6�{U���Bڒ�o�����LF2�
M]a�'����Ů@��XD��+3%�4e����_����2�yȬ���@)!ӣ(,��Zj���\]�9�"J�;G��E��5L�_�x�e�5M����<��ORj�c�å�M)^ �۠of�vik���l�-�h�¦�q�wC�jr��4�PW���h���]
�;���,���vG�@��4ڸR�rɃ�V��h)��A$�1���������"6���ӿ�ag�K����2y�Z���{�(�]7<M	Z
��A�#��8.q��9��SԘD2��Z>'�d��A�a4C��j�x[�@X�ۢU>�m}n��4�ؽ�:_�cD�*:�B�
�����~ڵ��ȴ���$`8���V_��<_ ��6' ʫEiO{�(#�6$��詩�^GjA�K4e��)�i��^��a'J�dN~��z�쵥C��4`���<l�v�$n/� �� �41�R�-K���%�o���Py�d&��O��l��
��YO�%>�2��f�l��E�>ü��q���Չ�cb:V��=$�>i���t/=+�	}��'�*�7�^��Kڎ��<�&�~����]`�7���"WNx~�� ^�)<4�Pwb"�<�a���R��Tc��ܫ��3��vw
�M���.]VU8�񐩡f�,����n�vH�̗p��Z���+������c��G�u��N�|�kv���@GQ��}+�"|m��&M㖬V焖��g�[8S�^��R�(9�8z�EGt5x�	Iņj�o��D���rcM��֠�M���D��g֧
��a�2��0����=?]����;C_��J5Ɵ�7��0T"�L������o�Ā��?��AW��bY���O�Y�l��^��ɜ�����5U�`o���!NO*����~�hd�PK�����%%g6,B�'>�
t<���qƗsh�h*��6���*��Mc��]TDdx���ϔ�{J�^�Z��}��pp��o>�M�Yi���z��S�����k���v�k������������G�j�w1�\����3`��+߇�K�Ns%1Vra=�p����
u��ԫ&�#P�ۣ\:g����m���!R D�l��@8��,�1ѕ.����������x��C��(��XP 8�؋t��*�U?�dv�����,�����y�]Y�*\r�y�Ϻ/Rg�'��4m+v��ɭ�"ɔ���(q����`*��#�����&'��1ʖ6��i��A���a����N�bM��c���G�����H=�e�b�G# 9K�qO�Rd�뤀�ў��]�΢@飀K�v��rgr�BN�ܲQ�F���lC�`�]�ʛ�D�V!� �8�t�����ͨC��&c>��O�dy�5�zj�&|��?��jZ�)
�����K¥� �1�;g�/�،�ؖ���K3�m1�t�23	 rt�7���!1UonD���K<^���һ^� �t�9P�Z�C�(�;�I$�}�*n:d����N��%}�7��Ȼ�缠���`G�\˪���~2~�����:��s�c��^VZ�RV���5h8�n �Օ<x�U���Yl�e�ϣ2�":NT�.m*3|�NȜU<�@,����Vl�9rcB�FN�UhW�ybE*��3A���.�j�)�/�E-�͵x�n�O�) >[��%���OB8�_+L��{S�������r m�տ#�]�v��ap�0��ƝH��z5��3�bW�g��U���Q���q@���*�W��#c��Ƽ�W�չ5�fϗk�0�2�6���������$��gM��\��V?[��ۜ>o6����:�w���g���s�BN����3*M�S?�����F/���8Jg0U��h�Wâ�fm��8�T0��6�V~,~
�C�hpHl�)Ȍa}�o`����`���6�)��ʥb��h�h�}p{h���t��@,�?8�6��z�0F�Շ]�gZʫ���F�Va�:��{]�|?����R��P��cr���pT���b��mա��FZ�4ii� ��Y���}#O=H;n
���ï�nJ]�F��#ѻ�w�)��$S=��F.b�h.��N��T�?�o�8�������z�4}�h��l)*���sȑ�Շ�}E^��G}��A�c8��),>�T[\���>�� }D�b��g��COf;�>1 ��n�%V�{����n{(s�1%ێ�|=���.D��E����¨ž���D(^]�ߍ#t��h�ބ�V'�ԫڀh���T�|a�^d}����Ύ�ͧNm��Gp��QP��K0��-װ@�TUB���9��B��h���v��]�)Ǩ�\N�J�E]���n��<v\+����(��:L3�փ\GN��b}����C�C��V�������l���S�s�?:ݦ_1�8,������Ʀ��UV����O���!��[�
���{c;̏��9�u�ýcw���fa�jt{>۹:�[���!�e��2����Z�tR<�s�X� ��n-Yn�B�v�w���:Z�`�S�i�9]bc��`у�{������!#��J��X�ez���wI9�U����kZeq|j����[o�M1��[k�Ԫ���-���0���@"aA�qF`��$�a��aL:����o\��^�)�iI#��T���-��R]��Ϭ��ߎZ0�_+��Pc1��.����BsI>4񇽔I���Y�S w��2��@��K�8����$�W�~*Ǳ���Y
�Em�n���T�:P�4�Q�i �,�y�c�� �-H���)?���.YC���F��2�+�����5�)CXH���f��g@�Dk�8B�����;�� �v_y֤�~�̰h��"^zɴpT�M4ˡÇ���n����y���wn��fN�t%�����Z�H�ÐDTY��J�� �b�6���G��o� <f�����Qm����p_jYɟ���so�zpOOu!4
�����݈Z�ˮIt+����΁�����]�F�XC��*�,!�zY�3J� ��k��AS����W'i�sWV��gp7��%�j���6�x�zm�f�D�'�v�n���^�^�BX]�~+u���h4��/:)���]e��[,�ӣ-���V�!}��\�8�ٖ����9��Įm8��G~Y�E�F�ZnpD�L��	�u�>}q\��������Jx���ǿ(�R*ȹw�{�~��K&l�0�� �5�Y9�� ��E*����$�s��I�B�0)�j!�e��k��&�گ�=����9���G�>��G���c����q�е�PS�IgH��pG�1�=��!\v^�vR�xX�`��
B��@+����#�}��P�<{�'�sJh��21Ȇ�85�"Rd ��{�x^��!Yt��K^��a�ʔ�t�/��[`b,$ Y��h�n\\���oO��R�G4@vbn43��qś�(�?<���G��-x��W�u�k,�ܯ��2$	�"(AJ��غ�7)��MW��kxCHeeSx\E;g�.�*�}�$g����~�@��)j����;(ɱa��t���in�
/��I���D#��aL����LqCR�i���>``ŋ��iZ�Q	�Q��r�}�E�`IL��Jֽ2φ�����BC�m](b�
!m{k�n�����בb���F��!)�K��h�j�w�V��x�u�*(X�D���r�Z�e�x��?�R�Zɐ$���k+�n���) ��R�E`�S|_ѣ|S� ���{�*�N�0W�s!�?����u���d��X�އ��,��L�f<Z��^�ѤVYR���8��f>��s	[�p�ZAFP�����d��/��K�@��=�zل�x~;��>�t�5���E�u9��k�U��Wg��5LoD���+*������i~���aӌ#s'����kVl5�V I����=S���/[�e�ǜL�f�L��<~�3���4��'|<��W.?_3���0Ƚ��Dw��zϬ��?���G�\��3�*�6)��_Wǯ����h��Ė�~���nP�h�����犺�d��ݪ
Hjm�����b<�/Z�T�>�*�����"7�����`��B��o�pE��7'���1��H��ݸ��	�ԇ����D����~�޾�����@�&��IS����󺩳�ż��K{�Ɠ_�H�v��Y3/�FF���#5G�k/�A$�!E�O֪*��):G��mGv�ɾ��pN5�����!����)H�.��
$[�h�x
 ���5�7m�bZ�z�jf5"+��s�j�i� D����솫��*)ĦXq��=�5p4�w�Eǡ�-�����u�"o��m-�۱9x��n3�0m`b�l��?	�k`?NA2����Q�Ft>�fDH;����HU G����3Mp���E�9�pcKn�s�!�!��aZG�Wo�������(�_�t�T
�N!^�x���5/�����p��f.���>m%)/���t��Q��]һ��eS"�l7�<�?�7�w�F�)�U�x��Fm��<=�>V7EZxY	_Z���$p��	V�Hr�c�!�S�����ٻ�GZbv�l.qv����;�(����g��Q�q�ȋ��(<�-�e�NߣG�����Z���U%�g���h������ө$�@߸滔!��oF�������IN3�����|�	 :�	��r;ἰ��J�r˪-��4�����HQɞq�_?���?��GT�%�<��N�nS-��ɹh3�ɿ��gg���TH֢�.�L�5�ߐ� �D%T�p�ڼ���C��A��Oԙ�XgX��a�X8�:/ '�y��~ ����"�Ⱥ�������T��@ʆ�3�uQ�.0�<]aѡ"\P��-c���� 6Ӹ'ɒ��ԇ)c�#�'��4L���ul�yJA��@����"��d���fė�����^zԑ�3�f�v�,��c��L������-���L@�U��?�*Ђ������ܕ?_��{kwZ[X�rf�2#�v :�Ak�"���l���S�S(L�AR
>M(��r�M����L�d��\���޹Xx}2����?��ٯ��XÈ:�ͼ6l��`�
7��FMƿq�.��KCoyZ˿����W�.�q����|T�zP�>C��d�I���
B6�i��':C�YKJY9�r�<b�R��R)�i����
�*L����lQ�-�\�`�]g��a�kePN��sg��e=�pK��;���S�R�a���_��,�]�9�� >l���i��ņ Zx>B;V�;k�	�6����;��L��r� �|P+���*+���UVk���������F�:0$��쇧Ob!�����y2_l\�j�Yh��G��tK3��WW+�=�*�R ۡ=	�|qJp�e�}�����ñ�k0�M����g���n��G`r!xƾ)��,����Ԁ�C���#Ӵ�K�o���@+����D6X��l����k\���`0m*}��a%�a~�Դ���Lg��C��E$���ҍ�݌��Un(�J���*���mYdq��C��}kuN�s�oj����F�U%"��<�4��)��m.`��6�M�VF	��EwC ���%�Qi�\�T��5���~�L5A'lºtʣ�/i�WX�L�Q��K83�p�O,q8��d(\Y������NR�2�=.7�|�
=�XԎs[.s�
`K���,��������f*3Z�Tl\@��t��[+Jz>;@E#:EH��C)k�(���B���R_G�W���|�:�׬~F�l�s�@Zo����{�&v_�<��L`*!���՞B&�T�nX�a���T��{�e��S/䳂{�ׄ���2�/������gF�=�B)����~�0f��T�#�}go���.�g����d���ί���Fc���<��JT�万�j��V"ǻ4��f�����Z�\I�Q�Y�_���ʋ�j<�bc��ch��m�l���V��A�� � ko�Kl�5��Oи�� �+k���Y��������w���cԍsr��l� ^�=6%��� {T�fZ��A�9��=�}ݛ~F(�T��S){{\.Wbl�Q���g�fࡻ�ܑ����ΰɛ
<����y�{����k�m8dǍYd�.��3N�t.�z����4�1��z�р�$����IK�x0�yQ�M����6cq�\˃����ImHP��Ԑ��<�I�/H�>���z��eH��pdck�u:�o�_�6�L��9�"d�Ͼ*B_{�g��9DQ4-c�x3���Q�:dG�w��r����#��|`�g�+���,3j��0{�2s� ˡNpC�W﫯��_9��c���*��N�⑳���`�z�w�j��U��VF����L����@
����J9�?�Ôa=p�(�p��{y��������,�tS_��}��gd���YP�/竭��	�~���鮻��܂��w��=�������W��@���`˙�����9%!	'�;����!�E�d�T�<��k�3�:�3����$`��Ύ08	ѷ�R]ٔ�sxx�V�Q��o)Wu~W4��y�OxH���ID=�������؎�ځ�����ٙ�+���N~��7$B4�v{�=k$:$o�� ��$�juq�A����
��pR��f����EbrO\ �
R�7�Pb�7!�����>�'���&4	�U�^���<���~����>;��d���.�[�w^�Y�XQ�����"�Y�G<�%*c�H��"�]��`��dUի��ؔ�L���5%�$
q!���sy̋aI�Y%���R2�xkh�b�<4kh~�-�k�!����OĜ ���5�e
�De8�$��@q����@�F�c�sX��`�fI&�d8��1=\3M��C�+PI�A��Dq�ҡȱ+�	*BN�s3h[9��6�jL��/EqIU��VRX��iU �:&��?ڝ�2&���K��6������2�T������l�gY4�yf��hhRv|7��$0�I��B�1��ģ6$��t~���=׽�\</Y���J��k
gh�~��*�ss@w&�y8A���T��8���M�KD��TYR��CUGzW�}�5xuۧ9�G�����G(V{���t�x�t��B��;?����8s�����Tx�e��kT@�?�Bp�nm�)�C�n�ļ��zR��N���=�8�>� ��O�&,|.k�q��djQ��'��2���]2.�Έ��ݘ�ɹ������+J獖A�&�G��1�U�]��ph��RuÇmN7��xY2���X 2���ks{��1Rk�k+;�ǯ���F�@�d=��s�yB�`]�~ȐX����X������>�Þ�e��j�WĒ({[(�FH�JҐ^<|aY�v�2��]�v%����_�%��-�ƃ]u�lq#p�{�|��9�	1>����a�f������ �1���e6�9#�x0�|j��,��7��0�"/��ֶ8�?y�~�ޭA����L_]�����q�}CKQ�Nbc�-��U!�h�WhMii⦏?cD�q�tv�ʍ+M�4�rfS,<�5��+��x$�3p���9���q��&*��*0j��L���s�������I����"|#����eQ�槮kך@Q�~�,�̂�k�M��h�a�� ��ig�g<{a~����!u��c �������F�f�e�&yˆ:Q�2/���?��k���I�0��$��9*�7�h4�܊[��C`fLH�j�} 3u�>���D���pEAL{�y�C����_rg���i׆��F���5�������M�TZ��o֥����zI�x��Y�Z�E��M���V�7$����:7�;'$J}����P�R9��@���5�v�̱�	���ނ���j�Q���]�Dt�D�b��D+��$��~���۝7�pI~ԩg7���Z���:P���B!�cg0��{�۫d���1g���5�u���Y�#����&�85ذC=� w`[h�)u6�i�A��O"aƞ���Ȥh�n:h �ُ�m�^�&ĳ)��(1�tת�˸�eT�	`�ҷ�����,��:����% 1 ZA![O"߅�I��u#�$m�z��U:m��Zó���)4��G��맋)Ȇ~AXh���@��]:%0G� @8'eW��9�p��s�Y]�m��r���\"Z�zyPUT��?ょ������t�2��+X�(E�W�.�����X����'=�ҕګFOr��z�*v�vJ�S-:݃�7C�B�D��Je �rU��ᶪ��BO�7RZnvFTd�I��i�;
�px���yFB����k�p%�#E�#�$`�}��\���O/�����Ugh�&��HX+���%l��Ro�ʺ�k�eT�V�7�*�Q���tO�D�~���w���xm9��GC���O���vv���M����[�y��8I��Hͣ�P�gq�Zk����� �a-g�'B�ܬp�_eQ7p�Uv��&���\ǙCK[������D7�~���Q���[����/��dS})ɮR�s��m3�=H��}��B�����?5�'E���	�ľ�dq��ʱL��$s�3+�ؕ����8>���H�{�@���w�a�u_0J��c�l��gU�2�5�^7.��B�o�&�&�tK��Ntą��A<���=��LӄP����2J-���e�~c��1b�P/����RD
Ү�E����'��l���[���L�EKe��Z>��i���o �[N��3�Ddn��߂��pq��R/z�0K�	%��Z��dܸ��W)��"�hZ�J��M�`g��u?f|ӣo�

3��h�?���Kn�i�S���y1	�2ETQ�������d.�+��әv\Z��Ox�Fte�9P��﬏ֻ({�-�%��j��7+��V3f�GDB6���4�5ʝ�<}d����T��>��������.b;�S��I��7�[��d����?�+�;�1���*�)�|��������{u�ҁٴ�#{쀺Kp�EE��DxEQM��PiU|�y���w��׭�������}�H�q�����1�U�T����d②n0���������$k&X�n��C����ّ���8�|Ɏ��,�^ڑ�C��N���ftZ�O^,z	�nF��z����IMô��>;�Xve��_�^�ցY$������e����
�������eK� B�(K{!�S<b`b��5ߨ�)F���� �I^Cғ��w '�g�匄�&�C�H�;��H��������F���� ꡎԩ1�
�К>��7�5�� !v!��Q5�N�=T��=��P�.�(o
��넻)h�T~-��3��/o}=ҁN�D]��"�j�Dl̟A*�el�S���b��m�*�~��H�X�V�v'L���	Mb��$e�o�lG/eﷳ(w����c���AؿN��$�LŪ.��k{6t�A+�M��{{���խs'��3�R�&RV�6z�8(�9����\0ʄq�:�!�4s�:[��U�LNo�	m�:�^d�$ƀz����F k1���(ƭZ�k.��'���fYu +q(��3���9E�r�88��v�9��վ�5R��6������C�?�T�o�#%s�PXn�zrX�w�rE*���T�1H!*hC�r�%�#�j� &�:�1�o�6Xk^�����K���L8ç�������Fm�0<���w��H�2��e*ݫ:/yN��?[h0H�Y�x��ݾ!R�-�<&���sq��?j��?=-���������=<��_�ℴ��-6P�Gخ���Y�U��Px��j���2�=�bUF����+�o�S+���L���5ر��6L`8��7��u�Y��92�a�e 
mI�ˌ2��y��g����u�ko��~��N ;M�8{7Ǘ�f�̥TۅV��S�=�����~Wm�~���5َ[��+�J�T�اu�
���^�~�g��3mJ+8����,l�fF�͆n|�\Yj�Uך�:�{��Q�n^h��|tsv/*f�ה[g$�I��6C��X/Nq�	���{��WJX��م�>Ѣ� ��t�i��lX�@�ٞ�~$�N�^^e���x��ITr������mY2Ͳ���4�a*��WL��"X��Է�n_��+�'�7J\`��@�e0,PJ5c0�Tœ���<@�gw^_f"ʧ� h=��Dl� Y���S2�r]�(X�̕T�-�E��u:h�������1�3G˜c-z���˘�֎������+�h3��P'~�́�����S@� �{X݌��
�����z=D:`F' �f�i}-#+R��k?�3����l�x��Gj�BT��>:��d��"���}9�����,�ԣ!dE]HsT��צ����/k�Zx��OSM{���Z�	�% \��>b(��fs@n�/}k�\ɢ~v���e�f�{�h���D����Bc`a��B���Cx$T)L�qY�r�d��.;imV>���4��>!. p ���iW�j0��<�xZ<�Vl���c�E�ӻbK�/���kl2�ݨ����6f��*0��~�������,�pK�0\��L���Y�5>���y󋁱J�!k���elm�䮅�w���A�������N�&�s��^=u8d'qd����JXh<L�O�V�`V��J()������Ip^� ��]g�[ҝ���g���f�"@EW�0�K�71�}yJ�9B�����77R�j{�"�<�]�$4��\���[
�/
��ôVWb�4�G�I��6��|��S*I�{�#��X'V_c�TO��mb��\��,�b�>�&Hw��Ɯ�9'@�~�Cԛ[[�a�UT��C�-���X�:o��U�ť�\O�~T�	�uhQ�X�eUsߙ�����"��^Q��= ��3=jS��Ϭ�%�����i|0��Կ��6�:�����5e��(�~	^�ZcI�%e��ک�"��R�N�{?(�dJ���p�܈��Z�4���n�mT��$�
���=�jk�!z�br������Bv]�Aǒh��N4��dT����J�q��[.S���~Z6v(�@�յ�~M�`@������zY�]<���p`>P�2�*�pN�C�
������4K.��coE_[��I�'޹lFe-��N����q�Ǿ��_Y�$6�����`�۩���/j�%�������nZ������pj�G���2�r�VFQ[��Ȫ������/�&���i4X*^$C���Z���;����a���C�)j7�Z'0�� �n��rO��o	�=`(�kw�7�މ9]��I-H��ܖ@}����v5kv��Қ�!�I�ZN��9�|%p�{��Xk��k�8�{ɩ}ق���b����$0��G��U�[iEL0����JQ��6���b=<5ֿ��
�O~����Yږ�#{c���5)]zqI����m�'��[:��"ݼ���}��0��ݙ��9��	�$�^�+�;�N;`�r�S{?��.>����i�M��gJ�����	�Y��Z��x	Fx�]&������7]�n�w�`H��f�4[���b4�DV�8��ҝ�EquH}d�>zra�ˁ2��7���5�-��G*�a����2�g�8�l[�CA��pܱ��s�x�4��"u�l{��'m��7�E�G�(��:����9��t�WiW?�Z<qV`{���L�G� �"�d�,TF��v������12v�G��`�S-5:Hg{Y+����/̆ͤ��<�`�K��ٽ�h��l)�'��#��Qۡ(�*�~3���>��R`n�c0��z��$C����J� � )�b��?~|����i&��wZY:�'"�����J���tKkp��DL�ʟ|VmM/^�)b��^I�~r:�!,�\�ǲ���G�'��ד��v6>y,W��Rn�U./xA�?���+{��1�NE����)�B9�{��ę7`x<U��^�� �t���5}�l��6>N�e��Ƕ�W�2���/�Yy�<��Ri+K"�d|����;U����@�WA����{k~ ��T�a�]Ҫ�}C@�:�>�S-Q�	�0A���UC��񲄟U���,�_M�ؔt��M)쩹L��J�a�2@X5qk�m�N�,�le-���X	���1#Ec���;lu�f�Y��EG
���ƻ�J����Pq�"C�<�����3�(�t�VN�Ã���Er�����<�����(��.�31���'�9�>$Y�R�0�g��6����m"7R)��7��Ft2\B����x�8�p4�8�����k�rP�ؿ�u{̚�� ̌�ae�����z�)��>5c[^g3lk'ekt��8)lU��j���"ÄG�J�q�|$>�ئ�a$$r��h9�kZ����@Ix�{��Qp��r��dC ��1�#s�dL�qѻ��_h3��!_XfR�)�=�i��QZ���<G��P�4O*ʗ�(o�|���l�:�!\:��e�1���R�S�@-hYN�Yȣj��_}HC��
�
`M\X�$Ƣ�q\��R�J���&^O���4��K-B6UN"�%�zH<DN �Zl4�9r��qԙ�J�y����PR<s	�s����3 ������*y����u�`�A8��3j��$Q�U
�`�����3١�3��z���\m� �܋
��j%��c�wsbAQ���Jt"a��p�v��$��7?����O�Q��ᘵJ��!�OA��2��$��~��P�Gfݒs���*�n˵���XL�]	����JW�C��rV�I���2�~C��,�hG�(�Q����A%��a����AhOx������T�m�����������	 /�����+��� �a{m[�$�d��EH5���c^��?�ǳ�[�,����X�^�æ)~ݧMW���J��D�!��B���/����(����2f]u�[�HN$Y�4nn4�t�u	�Jt�O&$,4;9g��֯*1ѱ�"�!b��Q5�Q��p)
S稓�2d>�b�h��ﶌ��^%�w�@i��f��i
� +��zb:��#e\q��91�b;K���F,ؗI���𣦦��$t���f�N��,��2R?$���R�����&�R��jb/�0��Ʌ�P�~�X����1��2�,��Lz���D�`Z@B�Z+��!��s���\&w�
,�w�V����2`\0!X���ho0-:_	����FĦOS�_��NN�(�w�ݠY�Q�'�7�2�Y¾qʿ��Ɵ��^JIR��A���Ѳ��Zi�iz��<}���99Ǳg����=��d\�tY!�|u��eq�N�*b_E��� ��~(�1"ܹ-�]z����Aw�l�]��x��~���|_!�P'��#/����HFA����������@=u��G��U��W�	���ۈ�^"���[�+w�?ȡa���͒@��V��g�	-�i��^0^�	~1H�D@��h��@_�u�rM�uᓊB=��q�ǂ���&�g:��ҿ6��w���5̑�@�qRv݁��m٠A�!�X3ޜ� 5�rE��%��L��K�B�K*s����C�gm�S%�y~ԩ�D$^��R��Gw���L�&0@:���� ���Rd��\2��-0H7%��������κ����،xjL��^:(��:2��q.Ta�=z���	���K�T���L��(WRߦ�h�#蠯�Ӳ��Q"
5 UeM��	�.&n::��&�]�p�E�^8c#0FFMɓ�-����7e㳤�#�c�����"`®���=���JI�xșN� ���(��ʠ<�N�ZXkn���P������њE�\����	oab��EJ�O#3�d����������OR��9>1��N���;mu�$��_Oի���Q˺��;�zیڋd�����.�&kP�����ꮈ	ƙ�bN�e��x���ڑ�o+��g�Fu(oH4L5ڞ�s��(�o����5��pM
S�,�[3)��� L�Z��⣛(Oy����f~���"�)�?��H;m�r�5�[�e�h��G�1&V�#�76��-��U��:Z�U�+�h�b���`�����Z�/�xlWi����~�lj�O�u\0ų_X���y���/*�{�F��f���Kh�	]���x���lt9��yY��0s:#�a!���mq�	\�ė�4ܿUI�:�BQ��Y�"�eK�ڇ���#^��<35�S�.�����Ј3��)�?�˜
U�L�?�G�йh[��U���,(c����	�f�y�A�Y6h8n���@��l6bK�]���V�¥�a��o�P���X}p
~�`���'�%/0��T'�!-���;\�O��M��tk6�J� �Tc�W�q]u�=+q�]�'��`*$�h�ٯ���5W�z��c���/6�Ck��e10�0|\	(  ��������!��.F�{�d;!��`�%�D���Z�ʬ>f�Զ;�T5�l�Q�M�+Ÿ�b�1e�1p�N��[,*c�d��p��-"���B�G �������]N�R���t�'��S�ơa�.��mt���ROC}aS�P<B>M�R$*10�WޱsL#z)4�ɂ�喙(?�&V ?�D71�I���Q�<��T�jX_�]�ӏ ��v�Wݸ�9 8�@C*��F]rrݛ���*>P�N�|���W�M\��k�=,��V�u��:M&�P���|�d�7uߐ�7	O�6K�st%�;�CTJ ��\ދ���Ŭbtv��Po������ʇm3�&7>���l������҇���|��s�q��.�V�9qp?bor�<]gi+�:�zks��EA���Cb�,bw*��f��j�mE,M+��]�*�n���W�x��^ϖ�t�V1�wM�&��T��p�bU��M�%̓KJ��Ά�]��˗��� ��.�>��Q�@��:q��[p���z�_��ʳ[Yzrp��
�tF���r��[�;a�)���v�@�`� �bJu@N*���z��F�hFd�"K_z{�/�W�r�	�\p3*�K&"���N��S����?�n��:�"�]1�du]�_ ��^�n�e����0�������.�jjK�ř�n�mn8Ba +�Z����GuB�M|��7s̱�Tn^��&���(��3�LK�)��;��F,!���s`��Q�hs���Rƀ ɮ}_7ߩ���C��O!q��.i�[|��$��z���i���D�e�*v�� ��ў�����0z�µ�%{X=rp/o�Űh	#�i9��~*����
�	g~:�$��
ر����0~��`��X�J�l1
V��QGX��k��OH+������K<��ǒef�ǈAaQ B��ʆ~�A�4�t��S3���c7s���h>+�t��U�#]����ԃU$��9�-�@���ݪz���zD7i��ؘ�`�0U-g7
=K�䜿�!;V��A\�?,�z��	a\�t�7���Mg�U�Ha�^ݚ�Cc�����}^u���4pw#�w;�$7��K�},�l1�!8��EX�ǴNYbJ̸�Ϩ�,-��ܥ��{ jIcD�:���L��D��� ��F\��e�_��}u�uu��v�D~_WwA�����y���9O��F�aҹv	��D��'�bQQ�������8���`��8��&���N�;�Bt�$h��۬��x�X��L�K��^C��Ρ�~nP���?AX7t���t6)��]ɧy����d���˘�8U������"L��ކ�I���ʊ'���"+���Ij����
̆�`�f�6��S�$��m�=Yjw~l�8�s�{�����(�f&函ɿ���1����	��b�a�^G�(V�� ��p�<��B�:�����x��P�Q%mi�d�l�O��4B�����z��4�0��@��2c�pQWøu��+/��\�>�a~�Q�XG-�&i�}�`]����|�=?�����5(�>,&�+HY= )sF��!6ڡ�k5�K�J�4M�6JW済�H��,�E�H̳^�\QmPI��R���2m� 5�N��M�U����PA5@�R�>K�^������l�$��`�3N��`�5�u��F=������MD<�v���&�}-�Q��6R_�a�P���o�y��Z�TK���[bK���w�zv;:�)��ª��En�s�Ã_��@��j$�H�G;k�H��P˙7¡Շ ��p<*�~�-k���}�2��.z����\�bH�7�|}�� r���jb�1�L4YM�e�e����Z|�[��}�	�����g��jg�\eal~�Nv�h�A}œ�ȁ���>c%/��=xz�Y)ң�Wvþ#����j�m��]{�{��2ű�GJ�<���ܢN��rN�
J� �&	̥����n�_�n(�(L�=sfc$> ]�t�76O�%�Z�ޛ�~l�Y��
�}�F�ro�!Q��!�<SHTk���Rg*D��2�8�=�!��+^.8�%�ܑ|w��{�'A�i��0<s"utƻ[|f��m�e�0�<L���(fj���Sj��	$u�1'2�"���o�����r\�4spu �;�;,��b�xs<��S9����Ӹ|���~k\-	I��VPe]���W,B�Țv��g��!7� X�W�A
�o�a��Q�!��Cpb�H���Ht�:@�Nl��8��{D�OY����@��H:x���!� ,�q$ё>t@րoi�F����n��B�]�b��~ ̯���n$9���cƴ�H�up�O�}fS�v���桾�����?ͧ�;M��w���q��P&�~��4��9Ty�;�c��ok�� rQm^�SAV!U���_�pa]:P4)���iZ�R�r�w�jB-�s�Ơ�=}�+��[�u��?���|4-_%G33%�)-B���	Y���|Gβ�g��y"�c\���8O��J�Q�¹��㳞屮��d̀b0��d1П������j�����X~t�:�4����q|Gk88���G%'O$}��zzm�]��ɵ/f�_���B�k���qp��c��3�sTɔ�Ʀ����_a�OE6����'~|��VQ=��w�����x��FW�]q�ju��d�T����	�7���x!AhY�Ej�2�ɳJq�:n�4�ۼ�]��U8�X~��1��I�������F��v��cg��;��3�t$���	����
��iX�/c��x�m����y�z�ka<�`�0�i`�lm1T��9	<dH1�	ֵ�ﮭY)�ɒ�ԘN[rS�|:&/�����/�:X,���Ii� ��!򎣒c&�8��=���6��a� �Zk�eأ$?7��1S�r��c���Rn cЌ�'yX�br�EÌ9�}�ɻv����P�����j�/D#�R/��$6�,o�L5���;��C޽�Ib���6'W�	��t
^*�.�n�2��
�n��EԓC��h���)ebP�:͌�x�I�!�Xu�Н�C����N�<�V��vf���)�� ��Z�mB� ��'����~�~3��V����+���|�\/��e��YA��1m���Tٔ�Z"F�Un��j�H���ke�&�2[D��67��f;�=j�\ ]���(�((4���v����(�&EiM)��=��#�j肫�N�C�7��v��a�$+�25�
.X4q�7������R�G8X �z�_���^�ί�<036�l�R��%:���j�9��W�	T+�p��ށJ_i��>�E��֒1�#��+�	�3�1� E՚��.�e-�Y�O���-.:FؚK��#�:hcL��T��	�s�|+����`��Iȭ�ֆ��;[�>c��ۚ��ޢ$��� \O�V���!Ѕ^��*Is�՗�@��L6�v!G}Ȋ�!pX�:T��W����誄Y��p��^��zN�k��̈]�M���O��4��H�DW�����J�P�M��z�������Z��1)���8ƴyx��8���� j8?��\{�@1|y�;��$��dr���j���@�i�����X�i�o١>Bv5|���Hī�O)ǂ"��p`�!^��q�>����]��gKu�t-�[��:�3o�m��զN���3�Ut�}֚5�J�r�	��Ocr@�"�E�����k�5F�~h�0��+�Շ0MaRF�kBj���V��	�C]5Đ�3Y�R�aE�k�/��� wd�Y*�u����כY����h��s�e,a��>���M�[�4a'A�a;��_㺠�x���5��X!l�J��^@`�4��-Y52ݍx3�F��X=��\��'VjfϤ����v��tφz{�;����b_X,ĊN�m�\HE������I5�s4�R��W%+�p�Z�,�-��}�؃���K8�a-�\����	J�ML,��a,��]5\K ��+�r��;�c}�~/��a|���PA��/c,{8��A�R0�ǚA�"܂V��u�~�X���W�\����-�<,� ��G*\��=�<�(0)g�b:��$�bg��M�����&�m��b5�m�Bܩe��6�S�+$����d��2i�*���)މe)����*@�U6-�4?a:	�*W;m$����?`^��s~HQ=J��S%��*2�R�_λn����H���H��}�7tt�~�i���	��Ԋ�x�}t�&���ft����%����U:l(Ӽ��)�ݹ�����-��l"�P@�?��H+��'�A�y�1�6��2���$RDֹ7��k:�Q��Gl�����ô��N?�*K����N��FN@��QDf��1
ێ�
��ZR�{�e*���e�r/��/ڣ����+��F2���W���'�~w΍9f��a	� =Y'�+#�`�d��b�F����__m87�Y������F��c+2N4"@��M�T������\#�{9oկ���gsޯ0��is�1�b����~4^�"9i�|G�}��� *б��s��b/P ��FK��Tl��'2Р���!J Z�ñ�ρu��\}�ӿJla%�l�����|�?����J�/�K��sJ�T��dMA��! �����t�:�!ꢩ��[&O��=�C���\.��)X���=�V���.U~����@�S��V���x>��~�_{���XA>s�F�_o�@��Z�����~|��M���T&�:�[DX���`�xȕNE��4hj�4�E��/�F�={:Y� n�TX⅊$�(wTyRZ���'�*�A�X��a[Ͻ���5[�8T:%I�5��I3�"$�|�u᡼9;��Q�poD��f9K^��-�
3y򛙓.�˅��ґ�	�ٳ MS��@�3_�<Cp���Aɍ��I�Һ�pn<b�aG��	�D{.>�aB�O��E_կ�ՙj���:��J�*�.�3��I�-	Z�W�1�l*��z��B��ǉp襒?�A�����j����Q��6l�������cl!;���oq�i�2��1h�2ԏz�l������X7�.wk�9�bWh�;�H0z��x+�")%֧J����I��v�1J�������:5tU���AZ�O9[���PS��t����1({yz�;��-"��0.��@�O�KIT�%�5�G�m֟,�G ��]:Ļ#;]u��i���"�4�/����v�F�$�Qj;(	�R'�'�cQ~�X���'o]�P��<�Y��V$��IƋ}Z����o��vI[���6eF� Q3XL!�g�������Fh��r�摦i k_�Xu�h�ma� /�/Z�R�h�x�x�z�����:��0{]��Ȓ\���ٹ�C����L�Ň�2�qT�Qq??��7��'����+U'딎�o� �r޼1d��
ݔ����ч��Ű�xF������u1�e��s�Z=���J��Z��9�YRd�e�{P�6�!q#���T��/�m�*��#g9N�T L����ְ��BRs�	�?��	�Y��=��GRn��E��G����gE&@��Z���g!6K��t���<{��N��M~�q��7�7@H��f���<�����.H�ȥm�<BО�"7\?��V���]���B3,��fu��{�St,RD�6\�u���h]SZ�^��̽y���g��� �M.����p�r��U���xs�����زG����4s>�Ѕ�WaE�̤�w��p��.�oe\)7�[>�9!����def�U�l����`������Z��8� _�m��o� )��]���D%����3�In@Z�Zٲ��Y����~�i�l��3�s�X��0���R!<�cǅ~�2lZA��	lL8�>߃V��N����l��K�&�����"�FB�\����y�Jćn���YӴ�����9��MM�os����f����_�v�����y�H�8�I��5��X�r&�ffy�:����I�A�������+�M����}2���R�*��c��<��<q�l��JeB��?��.�m�B�M�s�]:�^�_u]Dn/9�����A� �mh�{��V˻���LH�r~j1�J�H{�qPA��8�A�1���H�~>��:�}��z�9�A�� A,B�MX�A�Ό�U�N��l��3�[��ٖ����SĢky=n�-c���iYGyCp�,)p��o����W�Y�{���I�D��ԟ�@h��si2�W�.$氶����%�z�7Qm[�e��_:Qh��!o���8$�, ����｝S��D}?�+�E��EeC<���pV'8�R1�&�f��玜���zy�-2�/����Y� nhP�{X"���*��$O�_۾	�7�Qp��pQ�i(�� #���%���h�9��҇�j���l.���_��'v���x6M�������Ȓ<EUM�*�c�h����C�-������J
7[%֠)u�M��G@↯�~	d�v8�"��C��l���U���Q�g҈K�:������v0Q�\z�v�6��i���������`�k����n;�(w3�_C�"yY��e��
�1�s���	�X�9&B�(�{B��\>�d�l��{�0G�[���(ێi������:z�5V�H�A����l@'����R@h�=���-��Z�
X�������g��DLc����~�05 g�І[mh���YQX�L��5	�oƸ�D���Fig'{6SX<0�څ�TZ�'�UE�(�*\˨+ Sr^�N��,���;r�p1�x�0G�Y��`o�F|N�G �dvv/�Q��y79���B��dI9�~��%s�����D��E��F�k��4��/�9��`�2�pIzp7�i~,3V�Ϧ�65ˁ�P�f��^ 7��I��np�����l���4���<�oe1�6�ZLG�l����*<?GV^�܏��	�B*��R��VM�0^���
�S嘲��<�9<M��Pu�6�[�b�_Аh`6��^��Z��d�k����	n�?�8���®�QV� ��p�A��	����6v�5��k�)����꧸��y�RWI�(�;pl��J��JdiG��K�D��qS��f�V#��;�FA��%�jd��&�G��"��	y)�j�M���,d0;�e4�	wU)b&*a�h��*��i�A_��Ph�� ZU�Z���H���dP���˹"x�|>\b�۪�~ƿ��`�ˊ5�R��xeqZ�L�4#K�yԷ!X*=a��b��(�)�q����IG��х���2�'c�����e>{�����B�  � �s�u��;u�ůq�ɏ��\��'iZ尺��d��Ĥ�n39XP����f�!;�����ۚH��;���Q��ҕ�Ҟ�Ƃ#��d�>���R�9�&�j���P��=SM�:N;|�1�� Y�x��2gH�Jw׉#9B���-��?r��v﫹��Q����l��⏰�����t��Oh7T���wU3R�����~۟O\EU���^���!�h�qT��~��3d��^H�ǀ�H]���x�!��1Vt�,`1r�pS���5��M��$qA���x��<lz��P#k
#��g�	d<�(�X�4?*G�4�g5�i0<Ǵ�v�>O��9c�҄6���.y���0yB�7Q����M��?70y�{��Ď�鿵�њ�.mO�>������I��&����\����1nB��'=�z�����=nΌ/<����!b�c����j�)z����`�J$���p�/46a�������X�ʤR( ��x	f��a�*2#��7��&�35�.ˉ}_'S�^YL����M�$ NO�?'�}��eO^'�e]�ic�DBe����㗸i^��#/�����0 ���21�]���Q�j��-G���bK�w�n���V���KX�5E�`�G?ϒ���`t8��\K�o,�:��W$^Y��{�g|��2����x\V�*�C�8����㮘�$�2�栗*1@���V�"��ݚ�/9�A�)�����f��{��5��Ny�D���>�Sժ���DQA}�2LBN���71V��\���o����3[Y}�@)�� ��}T���fK�ވ��IEUE�o�mE�=o��I�7��N�z�$r���jR��m;I�P�/I�$!�I}  ap_��O6�G��x�7�F�&	�lz��E����(��ȜO����EL�[hi�SLr�-�]>0�%Y��<P�'���mlg3�vܯ�f�\M������2��{pWcϞ�|ó�C��x-����u�̝�0[�?�,A�2�^�X�p��lY��LL��r���x��6��Ֆ���ts�{L�d�!R)fl6�0*�2sfn��mZp%9 �R���G�M �n#�M���x����:��fl|��-M[���J�D�PJ�� �R�\;P�0�߃�B-~�9��mir{�.%d:��\�M3We�ث�2���jp�z>��QiR���hw���Ft������H���0�"+nB�$�v�d��Z�Smyq���޹��ئς	�%n��'�a!B��FshZt��+��7)�q�����U�엾:z/%F� �J�XG�Sʾ䥢�S�
����V�G�j�UX��ӷol�/�;Gh">��u2t�j#H�qGv�׮��':�'Y0v�CB�r5n�^��9L,.�	W���3���L�Gc�=h�v�a�j���r�F喣F����W�~�=���T�&3�Br����0\���װ�J�"�^���tq)�j�W����[0G]~6�]@J1�<����!l��(&��W&�҉+�8@�4�IB����3�k�m�`��Y%�1y��=����:��?ϩ7�.����ad��DN�Cd�<���?$�a�48G|�C^�w����
�QuaQ��2^}v�����$��H6KB����xdc.�LˢX)�V�$�N��
�[�t��)"Gf���myG���LC1���T�-n详�p�U(�z6��"�[�	��Hh��0�u#� ���b�KU�!����3-�N`����>�sJ
~y3�{2���f;�5Es}oL6>警��j��J!�n��wm����0����6���vv��?h�Z��z;*D��,yuĹ�U��=�m�:���!ZDH~�y�[B^!cZDnz �i�Fًe ���|y��pE[��A��]C������5�,�,�:�E���������|�V5�1�kK�������A��30^�@"�c�߳���W�	K�.L,�e�/�4�i6�Zĸ'��˹}K[����}o+X�,�щ�M���}���4�F.P�7��(�~�����'za'`
�iu����Gi8h�i�.�r:躍a��}̣P{�qK�l6�0T�D��>Cg�j�=��z/0��[Ȳ���?$ui�g�n�=�c'�`��2>[��u|<~�k���e����5>|��{�%爧(�M�ϐ`3P?�5��҉1a�����Hȡ��rG~�+qa��J���
���T��{u,�� G"�g��x�~�*�����Ͷ��e��y��{���b�c�"5�Xg���0Ȩ��wy�P��o��a�`n�~Uxwi�M�:t�V������)�Xk�s��t�\.$%���*� Rǽ6����y���Fr�Fv�K��(�U/nL���,D���/�&/G��b�J��esK��+ӄ��朧�P ����Pa����̀V�+ǽ���vv�o�Ƀ��={cL��V�#��g�2�ϑ4�wo���1�-&��O�����!�dm�1sԽy��	�x������Ykdap0Q�Z+
�OΙ����Y��ǳr�w4퇪w��e,eͣ|�s���@GJ����z��Z����dew�#T��(j�4e 2��R��H\���%���ʠR�ug� ���1��RC���+��?$Z\���n_;U�\w�{B�iP��pg������ĬM�fIR��Q�{��!�V�jTN�h���D�ao��0���m�'�k8��E��kvʃ��̚X����q�ɴ�꺥��>��7��8HY�����R���T���n�C8G���}�-B�g^��\��U��iì
I�3�][e����is��X����g�<�#��>i�ֺ�����
��QR¯�>=Vx�Fod���K�����X�����1�_Kl���ms�BSz�x���;M�4+�Vns������5���`�Bi�]*0�&s_.կv���K�p?ݨ�Z&� �D�T��a�䝑t��m���x[��[ ���gE��"�Q���^�ui���2҄0nH��eKx�B��9�v\:�b��?;�8��Z�@ )Β��|����8�j�����Np֠�Rw����1B%N����׳�;��6�/����s��D柪k� �u��5�"r縯�HjIk�!n�$��}��{,�F�+��G��Iq���/K��p1�!�{���b n'T��ƶ��x���UIA�46�cɂ�{��b��+�s ��ah��M>
�qzR���h2w�����F���#�8C�3�D���1������	�Q��{^���f�=�!��=��䎧S������E$)�!��&�=|1"ɷ��(�-�2��ܙ��N���/D�