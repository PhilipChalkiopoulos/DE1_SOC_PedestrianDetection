��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�)��7վ�n���=&%>P�!�M�L�6.�y�٬�w��5�[�ʩ�"��w=�e<�K�瑜�m�����F���М���dK^l]��+9P��D�]n�J�!��_�-0d�u�F:xY�y�jᣪ��]_�*r���ŕ�՝�U# ���G���|�����d�Y�e�>0u�Ɣ���G�W#���[n(�lV�ƕ���	�l6������S�?5RKj����;��]Z!�����B�w�����X�:�q�|��sT+��Tgf��SD�l���.x��0)ٛ��:�*�I�9�+ڶY'4Wz����Q��L'�������"X%�Wq�92�<�~�{�B_ �f:c*nn��{6I@Ñ�����������3قO�
�\�S�I��3���bk-`�ࠋ�w{�ҍ�_�5�,��̘�w�T�!��b����(�r�5$�Hid��c�|F���D��9��3��Ohf�<|���	�K&��8~�E��Il�v;�9"q�Y��h����p�s���ZX�c�tܚi�'�R���O?��T��m>���<8ᨦy��XKT�Q��%nu�O�k��>�<k�4�ؕ��/Zɠ���T�f�>w�-��d��Zv�o�#yʡ^q�Q`����@�'���4}a&���D;�#���=�V�b��P����}E"���w�˱�4���<���!�~R%�A�3_�0l�����.��n#�w�c!g<��N��٬�s�%�	�gdck<o=`2��c�o�z�am#�n:��D�u�~�Ò�sK�Kd�b�P(\�]*�g}[�kԵf>��mfҁ���8h��s��2�Fq��,���~æ��j�A�+^��m`��6zM��<zw�V��^��.�O_�������_�*�'�	�7���׈n#�n��O��,5$�a�,�wa�]�٫S�D��Z:*ǖ�o�qj�����SU�v����E��&��)p�ky>v��u%��{ʺĺ�T�.����N���?M>�)4x��sVs���+�F�g)�;�/)�Z��߱y˗�����������{X�{v��]R�5�N���ċ7aw��o[_��t��!���	U,;�>�@yfqm��c@��2ct�z�'���b`w���z�HW�h�hOڝ'�4���\s���:N*0�[	ߠ𕕘w�e�s6m���ּ�'4��F��j�k�3��%��єR���є��YYά����?�BH���M|�~z�9y'�"���D��3�r%��0l�_��0c��#$,���H~��v�/���P+	����z��Rx��F3��!a1���q�������cy�'n�E������+�4�-;�uF�g����*�>>)���dX��+��)�m��P���{��ډ.V�R�d&����F�Lhҋ��L�t"�w�6�@�1�^�!��.	٭]��*�*�%�$��;�|n�3�ߩ��L0��B� A���%1������ٗ怄 ]����Т4�R�o�ί��ՙz�%�Ӌ��>��K��E�T��d�+o��_�^�ǽ�����qx��س�7�6IeH_�X-F{pI���7�V��uR�����S�r{��������L�Ǝo��C�RB}�p�Q�^�%�b���Q�OXޖ��35���M���Ww��O�ks<�):�b�V3�J��ԦUsK�0��k����P�
� 1�{���Ah�Փ*�,e��ۚ���f4�Ć�7���d��<ƻ��&�|A��3W���u�*��~3$U�k�����gY�iz��������\lUG�$B�>I4��$8#�j
�݁ƅh]ؤ.1���/��ݶ��f ����+I�{�G�R/O?l�峮�G{D���	����hc����B �O�>Y��B��
.�a�fӂ�<Uq��'��@��������r�����T�*]g�jc������]�GWkq� &*�z�=�0�,ؒ[$񻋺�T�б���������������bƝWr��U-�H`~Ƴ��IJ��Y��xG�q��!B��ʦ]g�o�\<����{*�E�sX1^m��]�����o�}ѿ��+0q�f!IЕ����1訠Yh��F�^Q.�3ğ���<]z�(|h��fecV.�u��Pډ������r�h��_]�y�38�35$F��W�n��et��E�$��l4� 6���WZ���IÞ8��B1SZ�XO3���,��' ��xݱ��m�I�s5zئ�[1o1U���;��X��Jv�೤�t�N5A�l�s~�\��v�։3�v��p���¦���y�34���G��i~Kw'�-��%:m=]i���׻��Z��!��3-���,߰@�L�U�
��UvZ&o�̄�������*o;ǡsN7���-5r��}�#�Rr
�N=,g����X���A0ٌ�4e�P?s�{El,���fH���t����J�i
���^q�%��7��k�I�>��m�G@U�k�K[�(B;�7�U�D
��F[`Ŏ���F����i��@f����˝D��ij�������ꭣ�Lv E(�*������`��tP*�|CɄ�ju��e�W��OO�/�+9�z�?-u��8���FD`j��,�n�č�U�ְ���>OH��qGKwqo$QW�:�����4��1��k�aT�s(��m��.�#A�N2��@.��>�t��ةOmD�F�i���ʷU��������d� �-t���Ph�ȇJ�+��1�*�e�usjB<��3!F��ڔ�{����e���w�m�ʑ�=]�<�[��"�,���>K<�=��N��8�P�1
����/��"�>�,V].��쑪}.�����vh��X2���$�)[�Jo��;�Z�k��|?�l���� <�m��Y�J�L%���'�ҀQ���k_7��[���ʧ�
�v�g�֍ߣ���C���D��,)�̞��:׏S̭��w"nF�O�ͺ�**T9���#vz	����n8>�#l�#�L���hk_�Q��}�F�՝a�,���<`���J`3�}�;�ۨA���ji����Uu=�z�Q�%��i�����kM$��⒎�9�e�A�}|�5������Eu�p��)T�16'��C(��G�q���y&	�j�K[���{����� ��O^mT�֫b���J���}b��PB���5N���=��� �fď���.��A�:��R�+0��{q���_�+R�g��U�nB,K�1+����ѣ�k���Ŋ���2&'I`-M�5I}�r�C�i�put$!��gDO�-�6К���I�	[Xd�~��8�j��Rj cZXTvd�J1d���X|�7(�:�巾�O��ŝ��u������[�6�����)l�I����[>%���Gc�d��2YR�?�J7V���p֭/_s��`B� ;�p&����Yn7�,Lb©m��&M2Ab�m页bcU=-�:B�Ľ���k�| D��1U8͟�t\u$�t��Ü�Cn�EƚU�[;WH�:B�JG�Q�;|��|���J	,i�T߸,#��Hט�C��;�i��78Kֱ�@�O�p��>߄A����ln���J�ew�����;(M}g��"D�^���	!H��"]�ض鸕�xQj����:)������1{�=�~�}˟��H� �Nʿ�����"����#�����P���,�HjT�˅����,R��3/��:x��]f�	����n��ì����@�|�2�ֳ���YK;��@E�l�i�@D�z�&�M8�ĭ
��o��ɺ�����X�FH�~�W�Zȋ@�8nz55��W,�4�Ҡ�v��}��S�)q��=Ш{O���z��Q1dĮ�z�U�ޯ��e�"�fBK�ܵ �^��xZϕ3�E��t��V�5�j��k��l旵H�e2<'���C�����k�嬚�`3��D�2��]�_�.旓>ho�s���y�ԤX�'��8�k2����Y���?W%yM<wFNfV��r7�4�+8�!��8�H��.C-H�=)��W8�O�L����Mn�ܾ��i{� ~C�Qh�į�K�ɯ[<��Q�>�5K�`���12	��ij�,�H˜�WY�E�����*��95*q���:Ygloȥ��H"o������N'Һ��n#��17�eے�A���{S�$a ���]{#֎;	����Q�b�a$������fe$9��+�-���H ��B5�59^MZ���E _{����I�EI'd`)t��8=�É��^��A���6���s��p�AS׹7�EQ�>���\3��>	y�ep�bv~����r�������7Ja�����8��2�da��d�+������%LH�@Û��]v��ġ��B���m�ǎ��m ����f�&ϲ 2�]ݎ����h�
M�TeO�s�i?82�s��Y�Ş��w��ٙ��4HB-S�f���Dp>cM�%��F��J���.=�B�B^�_�O�gFd|��gt��2��A�|je�À���0��WK8k���Ů	�>��W�sb�$�Mm.>ٲp��@�h_sr2ֵ.J
��s���2�R���"h��P��a>�:ş#;w&������Z�0�� j 䐡��7��}�;�$��q'�-e�,:����
�J��<o˓~���ڝ���&���E�аf_��.6݂1�͞�iCj�C�3@D"e$���oD߳�c�ZW)ݮ�e�8_ܳ��f��&�qӸ�y�3Ug�3�W:�\ј���Xvq�c�8�>,`��>��s