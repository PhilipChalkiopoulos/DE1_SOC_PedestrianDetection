��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X������r��#@�/�����4�p5���4;Od��N��r�I#��7h��$�(��?�g:�ZGY�bӍ��0Yzb0o �Β��A���p�6� �����4���e��Ǟ�H� �a�C���t.����+^���}��G�|lm�.�|����"��(�cx�m1�#�N�N�:k?n~Sn`�'|���y1/)�
x@���n�+J�\O{&	�.�B䛄�%��i�f�f�L�u��i/���R�@;C�!�M*.ɪ ��_�zG�ȍ��ڸA�9[Íp���="N�jZ��|݈��y�A���_�������ⳤ\B�ҥL������x%��}�D��c��t�s����PF`�t|����Nl��W�`f2�C3�$�IF��<�Χ�[���jY9 �$Rv3�4H�6\�&�;����P���f����_��r{�M��-
���Q�V_U��	��@��;�x���!	G��Cm5��F5�Xn۾��ˑ�'3+�����#��!M�v�Sr��_AW�b��I#J�
�.��l6pJ��[��[���)<�ª��W�~R�T�F��=.����f���4���|��=W!�kp��T��Ӈ/q0��+���G7"xX��6w�	 ~�
�aǽ���?pŇV���e}ko�X)2�y�Q-t ��^�fOM��w�V��tO��.{JƗQ�]P�6w���w�o6�U��u@�Œ*^�8���ƚ��v�e��f�<<���7m�11��<�Y��ԓ�����8�20�ΠVafC���ݢUK��*��z������D\�yf�Nb�������`�ȖD�I�2�{�1S�J;b�d%`Z�[��G�*���#��[����i�CKA�
�wy�7��?4�vAqN��\
` ��ɍ0pV��r�\��3T�(���Vk��fo���b�-�[͐"b�>8�>`!4:\*j�����r&Es�� Ύ* 4T%6���;��FM�~��z��bd�)�iU:rf��HҼk���U�w�Gl&eD�x�=����H�jK{��4m��Gx��U��	,��I����`�v����F�t����m��вUH���LK=z�G~��;���ǙtG��n1�CoFc�w/��!����%#�~���P������\1 [�&Ӎ�v.yU��M2U���m3U�֫=�06P�<�j%��IО0� {wN�����s�k���7�*��U�]�Ty���~�-{����Ԫ��a9�@�����U���8]w���$��x������W� yY��P<\B�V@���"h���ف:T#��`������ ~�w�,�5�1��y�+�g(� lHwԑ�(G���{fu��~�����k����mu���:��|���Ӏ�H�P�(G<��"G5uW=���m�!,$Guߴ�~�|�D��#{e���+Q@�7#X�A#�����Q%����/��b��J�O�F}��gj��������B��|q��%!��z�$Ivk&����+?e����,��(����v_�`�*�Buȧ���9CL�5�r��g%�~�ѱ�Xj���ԧa�ƿIX��G� �D��h��^;+�8��{4��#		���n�j9Y��JE&��VPJ�����#��7.��Z�j���u����a�����?И� Wo�?��S�$�w�������E�$���i��]zk����1rV�qv�'�隷l�g�]�86Od"���},%;�J�C��>	&���YJ�)sł�4����pH�0��<��Oq��|"ǋ�)b�<?��XEL��\Ȅ!��Wi��p~h��B����z�q�8�E q��G�� \�V�ta�p���b5t؜���Sa��'��׎s��<��՗�
�З�#u��I��\���9�y#.��@Ppk����|�r5w�_r��݅�n�ъv�Y�?&�O�'L�>V�6��Q�`O�Bg�a�%��mEc{�9��d��gT�b[�p8�5k�ep�iLLFW�Ƣ V��՟kAሤL:�GD�f�n��ͣn�
�¸B����S��/�6��	U�Uڱն-Ge�ǹ���[)��cT|�����W�������>� ��x%��qCI3 wT�Y�|Rp�R�dE�.1�rK�0l�>{�B�(�,/�3��+��R���a
���FYC�3@(�`�z��x���"\�<Rb:�h(!���8l_�֚g��|�CZ���Ҝ��j��o�>Ƅ�X��I���ؿ�$,'a)!z�����n�u�e6�S.�[��5MtmW�cI���^ ?�<VQ�1�@W*�YM^���ۑ����e!�^��6D?�������u~O��,�|F=&������}տS��sD��G*Vv�ѩr�����!�kr�V5�-��?�z��TU@}a|��W�4�͛]2��*����cb8(�@Һ��.����[���O�R>�8�z��l�������AbKiFU>���wݏOq-_��#�4�2yQ�~.*D'���4���g��v�RJ�������7�}YY	V��T��"��QةwTA�{R5k���K_�`�$>=�Mlڑ⡞Ә�U�0;غ�_7ЧSUi�8J1klT�;~g���wIA�K=R&u�UͰV�x祀E�%`<vo�!�ܭ6	�@�7��/���l��)�T|�Er�7.�
‹�� IF�����q����W��.ͮ^�D�	v��:�B7R�@�BE��@	V�0u��s�Q_g$���^+�N/)�5����)M�xgN���sҁ�qk�^��9�"5��U=iSC���|6j�
6ax9�J����_l��
Q�'�4�l�-g�#$�{�W0�NZ��A��R�b)z�.sm��w�K�����mi�O '�T/��V��p,�ڡ�]��Hg�m�:4�~���&�ǯ6��OL93W'�2�~��{�d��(	��"�������3�������}˳CuEZ�ثI)�P	��=hxVKBD`=�KL��5�I'�e�<�&|��r�w��|ן��A�+����4��P�j�شC�.�D"��|�k�`����|5������c�٪쳻q�|q��B�?�:��)�O�3Ј���~q�����ǣ�R`�:���	���Yz�ǈ�#9 f��,�]8'j������!�l�$q\A��+�׏R����׸	/9���x�V�`2*_�D��k�����џ���Quū+M�ې��\�zm^�.��K���&�txd���r˩�S�~�p�]y��yCp�n ���<��뀐�B�:Ze]�LI�;&f�gE��5��?�L� b��?�!�^����k$[�R~�L����{����^�4�7c������I�5�-���&K ���֎�	�+��^g�^�R
����])p�BE����?#܉C�\5��CW/�I��=��O�zE���*q�3R�䷦��u�Jz+�=d�f��d)A��@%.��Ϣ@�>߬2���:�7����#SN�U�?�ڲ��������L�8��A�����f��
)����I�}����(l��k���^C��*�9��4���S�^=�wꭍO�l�؝/2���<m�!� dܝ�m^�8�[�:��<F?D�0qq��\�U����bV�'�z���?�Y�N��l�	̀2��3i�C;���3����|}$Dh��^��?X�6v\�C��6���Q] D�A)�	6Q�\��'�~<R��G��'1�C*߮z5@'LH�ז���қ@�+Sq��?��ɸ�R�3�f HL�"��*%N(��&>:��ͷ�m>���:)ܗh�iΪv�&��-�s������Vo3�>Ż�c��Ig�����x|
�fϜ���4�����D��f��3}C�}Q}�a�D�O��k-��(�!�퀲�����Q$�YH��P=�4�%�P&@a�	���ipđF@�<�ϳ����D�9WZ�'��S�e��z���^V��Ug��2l���O�֦������� 6� ތ�f�-�R����j-?r��	�j�u�~&e���-�������k��F�(Wq�nފFD�zU�W4��C ��15-SM�5S�e���[�#�kש�`�$H�z�3,����~p�6�Br�;��d��R����h	���[���=�Nd2ΐ*�_6��4c�s�$#җ����22�f?�5�1I��L��p��޳L���ȯ>�-�"�����)3�}Ǝ�Ш[׏<ց]�?�r^&BCbn)@;��3�r�\~��P�C���Wn�-�ݤ�V���+�I�3/��szup�䵾1������$C�	PǦ}������a�� w���`y�%Q{��3���ո�BXݲ��k���3b~GV�0�.i�DT~]>��Z�"1��I�h�d#�~����Hx[{(�:~���JLw?��EIЀ�P�ӷ��H�����S�~�W�OVB��&^m���EI��Ya��v��ґY��t3:`~�MM��WvG��� ��ڄۂ��亵��LB��E�X+��L:�D��w� ^y���!]N���o�uw��j� �[�yv8�
9:�+�o	N���"q���b��݆���s�r�P�(C�}+�Ÿ	���c���=�M'%�(�+�=�"7em3��p�
�8�w'��*8�]}�go>+n�s��@�a�R����xyQ��=i��t��������H�xw�����n�+����TQS�>�|*C�D��{N[��f|1����2�E��@�W/�koA��{�h��ΞR�W���n��z����lg��Q���A��H�v�V����+`L���^�0�頻�w[�jRJ�p�R��@�;�.p�VQ�{`K���6nS��0��c��]aA���Z��s I�ϖh��.��q��[y�9���ۑ�U�<�_X���� 7R�� ǂ�	�|�4s�t��Jd��ׄ�2W�Z��983tu��c�%���9�^&��PY��0bW�>*9�3�ny`e��t>�s ��g?yPF��WL�5Mc@{�3��oX���9�wA���}���>�P~���y��w���jhG&�-n�K�!]2�|�%�V���M�E�a�=��`�<U��
�\��	n���F������5��-�-��)W󩱉6l��[[��9E��Ts@�Wc�����K&��w9f���گ:s��*�*!����9<��.:a��t�>�G�nej"w����ue�g���2�ƀ�1����ϺE�	�R$���d&�V��{����ǂ+)T�k����ڈ��<�;��������汚��d�0&�pd��+�(i�����_�]/�ò���[��S�3����3�O(�#΢�ɏ���h=�ڢj���y��&�i~Z���8�Z۳�w����0+�d�s�n�6���'��k{jk���玧Ad��|�Q�\��5߫E��{�ܿ�F�������ż��\DV�sn��X�2�O��T�B����G=��uRx�R�E��c7���ٚ7�S��V���VaE�i+�v�2b���뀔c}����jWy^�?���9гZP<i{��]�7�xQ�K���C��ZZH�D�ϛ]���G�olO|{`����A�00%���L���:1�@���Eu=��v��%�??P^�m/��Ϣm�3!l/�3��@
��e��bL�v��$W��;�T �§�k� �W�]V���lq30�����7ϑ%[��~o����yhTe�$��u���zF�]L���Iw���8{h�h6T��-Ϛ�:e$���"C�U'�-��Ƕ�Y<^��Uv���}�O} Ĭ�$��?�U0��.�6���Y5�x�FH[���+8���m�˝�@����J�p50��k�ÙP��d$ƒH�&�Yp>�s���v�Ġ���&\A�Q��|��t��
���izF��&V:�}4͆�2qB�i�E��H�8̤r����t��N��fKh�4��W�T��$�������!Wlس�.�1��tu-`ADU�ڕ�Kq���p�~���di�����*���.*޸x�\ �_��[K��o[��"j���걕�Lڃ����A��r
����Ů�%J����Ӕه<4J����"��"3������Љ
iR��Dx��=��T	�\S���+��E�r<��XU��g�q �~�#���f�>jhw����<��V��7��Q��-�E�x����G�f+��T�j���f�Ǯ߂ӦA�65̟f^a��d������^�'>�oRMl��c�0i�e}�z���\���H:�@�Ű�bB�np�hk�V��H�M�7�v3�MT}���
Z�L��?�����"J$�y̚�R0_{͇�E��E�fF$/y3�Q���}P* ��#���R-#�߰�����	lT�"�%����&�$��Dn+�D}$�(oV��4H!��a`����c+!0��4V�E�)������J�3<w�I,OEk=�������aCW�ɢ�5�"�X�g�,����r�$=P3�Ha���A*p���8\]���gH�N|���d\� �H�X��6� /�/�\<(J!,/#d�ˑ�AX���/�v��z��Q>���N�<��"���>�"���$$t�J+G}�"�-�}���k^~��"���M���꒮�*ߑ�JzU`�R*
�]�������ۖ^�fIm_���p;�*&�C.lBe�R��ghDt���~{�qB|�;G�F�ՙ�6�
d���=-HW�\X�ҍ�������p�y5c��$j����j��0Φ�ƀ}�a�-A#��٭�:�wNӓ�x�~%��J��)�0Lm��
W��j.���9��P���Ȼih�Xl�dtS��8]7����템�i��<іk��T��C�ȓt3�j���<J	�7#�rߤ��>�$n���r�jvUӯ���:�p
�e��x��ك�����C,)��-c |�P>�Jlu����g�m/·ʘ�9��&G�&����o�.�hK�v4R�`��rU;�OEV	�ٻ�	���[�S/��S&˻�!����I��$^�������=CˋВ�Y�-��F�z:��\v����7��p����Bj�A����S�׶��<bF��wh�f1_��
^�?[G� 
{�j�L�`��+�ZjGʙ��6t��n'����N�>�e��]�B�r�'�<�����{��\2�(S� 9ab�� ��H�XioZ�Z�9i�����Z�I�r6 ���G�^O�dO&B��5�6� a�9�� �ݞ��¿�U�ܛ��A�dQkp��{s��&���5pK���v��"\�[�NdhE�[�Ȃ;R�!��y@H�C$'�}	�7���gG���
�9!�.-h.X�@�/��>C��L�I�K(�0���{����8å�طt����v�r��g��}�_,i�δ���߃�L:=�rZ%1�'���ևkm�i�y�,�2`%it$pnsy'�ژC��.�p{v�`*1�f�UD��\]`�J|ȃ��,�Q�C���� �\��b:�1!�"�ZV�O?�A��~��wwKo�nS�z�U��3�_G�>-�I@Q�D�?����׮�%�_�qQ�ë>/\%�P���w�Jlk��?!��-��`��C�q��JsYV�,�'h-1�[��0�:���	(��B����{k:��ڞ��4K�L�Sq����s9?��;8,�K������n��D�?�@�l
W�-O��?�Z��¹����w�Gn��Xz�oǜ(�R|��f���2u�l�]��®� ��a#�<�޻�UN�R[����A<ŷ5Rղ�̓�� 7:O9� ۻo��g�,��Q3޲�>M&�����ɢ ��i���G����&�=
c"W`}U@hk+DQ�8��K���{��͏�|���}P���x�J;�����~��*4�O��}3��A&��yJC��i�>U��;r{�cITP�����T'�jEFKRQ�(\�~gzsv�������Z���<ɻÆ�+���_X���d˳ҋ��ۥ���p������j����6�c�K�Q�{��0�3^��	�ZSTcSo��s� �e������q�ȹ����h��HhϥV��
�X$"S�T����ꢑ���1��G�NG��m��]���Ĕ{2��hD�>Ű��o�R�1�H<*��?�:�Ot�m����ʥ�9"8i��4�kC�n�b�����D���y�H����耹rnKu��*^0���aW	7"�
�n�x��J��C&f"7���Ph|6(���L��N��k��3s`�BZ���r�}3Ϲ	Hg�A��Z�$����I=����!\�j2�v�i`[����q����G���Y�~��� fvQ��m!�KD�QU,@����#��B�~�D�K���N�6a�`$�^]�U��6�kp��O��/0�=\���_�.��ԉ����`��h �r���qю͙|'�̉Z��zZ��,%���;�ܣ��>T���iܖ�Չ�I'j5�gywK1�ZYx��-"�O�]�9'/���(���4�<?�Gĺ�[�C�M% !7$�W�4p�1��D�3uz�S�72L�=˿����5^*)qGaR�-���t�R�H�t�J*i����g[\��]�k]����e�A�:>S����,L��wag_�}��5��d"�U	"th�\=��,�dճ�;���x����T���ے@�$M�>}_=�;~(�I�k��\�?��Ks4�He�U��G�� ٰ��jP&�h��gښ���n��刔���RWbi$%����t���TN�
Dj4�@a���<b=�'%Qw��8*�Qe+3��x�>Ԋ��lV����yѬOQ3[K�ͱ�e�|�zcE�c�\W8Z���������	��,��%E�ce*��A����a�_���d7���a���/��H�.�4����v�4���b$�զ�-�ի<8�ɓ�pAʸ���ƈ��9L�΢G�O`d)��z8	V-99�G@Y��Ryh&����</N4�ؤ#4ȯ �.��L�u�SW!C;+����[�C�}��@|��@@jW�o=ZW��`ت��#zP�:���nF�9s�yC���̵4�k.#�	��!e�Q��AK^��Μ��SXV��]�74u���~qNz��>t���_(/�B0��c�m�(�K�5�G/�����CưC.����E��'�5��5_06��^��͜꬙���8��m��	Hw�0����F~��Z���E���㴾DrTH'�a�%��$�!�S��Ƙ��7u.�L�c�/3�Z�Udc�俨(�ڰ�[�=f(@�$�V�&҃�M<���x� �'"�w����=}��iclcAj�f�H=̕�2:v#�5X�g��5�m��rg;��������ܗ���ƨku_>Q|�Mo�G�-��m8�)���2W��>�|Ngp�um�$#b��;���!���u+�&��I�Ȭ�*��2�(�?���H�~�X��ʷ �@��.<�Xm��<w�m�����g2l�A�zj@�hPUJ����͏V�X�Y݁��Qb�@"��7��-�y�������)ð��2���@��h�0��*�9
	��|��{>S�*�&���N �_�P2h~��<���]�"�?�]=ߍKܷ	Ue��|{	��^���l$�Q���F�7]b:�UD�䖳"!�����o� ,��ʦ�x�%vZ^y.�7�E�I�E��V�	 "U�~�6�O�
d u� b!#�����7Ƕ��X��Y;�=��Cc�Z�5o��`þ����4���}fp(%�JJ)�}�E����Dү���R�Y�+_=^�?�]�y7���`�V�b;��*>�W����7�)�>�{+���� �>������-`Z���R��	j���.�G���6�����g'�'$T�6�F���+08�y�	�+�ÙT�G�/�B�4�������ҭ�������`B�t#���� ������� 2��j�x�2R=��з[�[A�|ovS�0�PhɈ�����M+����i�@:�}�4J�4��"�_�s�@T��&��0O�G�[EC뽩��cV����㝕3�x��T�jnp�e�i�$;0���'n���M����V=���rE�e���o�����V��>��P���q
J�ʸ���r���o�)�7e�9%#��P��tE�b��gcF�͛lX��[�W'�5���u#R�	ԬQ���(�12,*�;�ÑR�3G�bQ'N R�F�T�G|�HR�#|Yj��bN��ց*�i���s�QY;yw�;` ��iGմ��v��`�c폠��u4|��*RjG�>Ԉ���Q���}y�5K��(��O��W�|.dֈ>A��e=0�\i7��O�xfj�	�q�0�җ��&q@l1�<�\�w���\b�vm�\�6#Js��0S-�t�bD�]�TD F�%-�JQe�1���8Z(�l�J��`�{$�3XT�&�v>�d�Wt�H5��G�ʫ3�5-xE��H�j�q�\YQzb$+(7,��BP��_Ⱥ���.����c�` ��r�U�`��ı�$'��g1V ao4
�Hڮ�U���Z5e1�WW��!V};�-��1�b����:�8�Im�\i n��T(��|�m���b��-����d'��,�R4�?��#g�EF���Ӛ�>Ts\'Lƞ������n�>0 @�1W�:P�P�$�6��*g7��Z�F��ZCI4lr����]��Mp��S7�H[�d�?�t]m�R��<p�V�9b�p���-\�hM�>੺`\gU0<�9l�)�d�L�ḁ��U�$�w�c���l�E�<RJtS��Y����KU%Q���+���Fז�R3^��b˹�i�zZJ
�O�-PD:@��<Rg�7P�.5��F�A��P���S��"�	��R�� �wt����s����n����3�kh_�T|��&ť��:�4�Е7&]���}ذ�xE��Nk�����]�E���H�?���� �K��ृ��2���=�v<�C;��#�xP�g=w�r K������q܏�'�����:�g��o����TϨzC�5d%��˛�S!qƥ��r��pe2�AsB��r��mb\E�uo"`J��K�x���)�&��9�P�n�t�9&R:��	��b��	�i	̲�C���!	��=ƨ���^��t��Qo���:��C풉�)�[��ZtB'���R���K�!�0�[-fB�ۆ�>8WS�曆J�����KMֲY,\���i��n2E1��JY�1��~q�R]�@�2ձM;\��&8������Y$�����+���}ް.BYj� �v��Y���oU	�bc��";G��c-t~��w�t����tb�d�@X2;���EgF/����l�˘��;�RЪΪ���-�<d}ݯ�x�V(wPƄ��كv_8(�/#Hw��g� �vN2h��	���U��=��Dw� C���a~�{�S�O�\E@��X>���X�������Z�2r�7�J�����ܖ��������tV��������v�M�T㥊+4��Gc��@�gD7@#�y�����Va�정A.�Ȭ���y����h[XB�����`�$��S�X�d��q�������Zm�� �\fZu�*�[��we�G�q�����JI(�*W��Z���Ɛ܄�WM<��_0u�e�Ep�����y:-)$%^��؂$;1�TQ��i�Rm%�O	3懝�-t,��;C�#��sEsf��OqC��Fx�Es������o�/ͳ����c)��%k���cQ�8˨�VE=o�������+`�$8���Bt@����|���p[z���JR
v�	c�gCY2/@�!�N����.��՟�����R7��^������sT�P�p���HٝaA���Ŋ��5�]�6�z�T��bP9b�Y�6gz�4����wC�ud�CM�퇔٦�f�<w�BUi|��o���%�C���t���*a�dWc'���5N@�Gw\yJ��_[�0Nx�?�p#j´�[�)�ArN!@)�F(��bҏ��;!�)PeA�]hĨ/��, [
\𔅴�-�P��� �d�Vt�lz�R�4��r���wp[U����ف�J7NNg0�]C�:B�#&���it*vh���P ��)n��K��#$�
��`�nz7�qxc��|U�"1T;J��j��{�K�#�[$��s�e�;�������Kh�i6D-Ĝ���K=Nj�q&U��Q��A�U����P�+X��:�1�2d��cj����h�RQo'�ٓ�O������%�t!Π���0Ds����u��:`��z�&`Ҽ�e�)��C�������OU*M�x��2���7]��4��(+�>�'�v�9��6��;�9�vK���"E ��������N���pS��!d@AOh-Q�i�nޕ�c��X��@�CtS��X���k�$)��d����Ÿ�舧آ�h"�0�����BЯ����U ^�P�s/��i�0�T��3��;�U~?-}���8�s,�������	��73�T27E
�Rt��I2{\yavx.����TG���k�Ѵ�Ϋ�~� �~��"}����]w�h�kb�wY��rݣ����;"��Wf%ILL����ֲuRo�˹�z��m��
eE�f%ý�Q=��Y;��^�������p����fY����n4��;4�5J����}쟴U�%%�{r=�?�M2
��	�($%W�~�_����4�t}/�S=|k�!��7V��2!���ĪNE17��{��%�%�x�y��	`q���b��xj�)�N���Ŀ�nD��D��`�����G�Ò�$�];�u�Zo�a���ي(�!r����\sSo�0��w�QC�K#1��B��#d�_�}�]F{��1^ӓ�%n�<��r�p��$G�����z����q��3�cn��Wln�Z�ˌA��e�{��Er\�Pr�s,����6Z�M�Q�γ?k��Bh��E�A����a�r����^���1`)��I��5vYוZ"/��C�,��"�7�f�6u���&x�֊���Rx"+�β>�xj���fp�8Q		jm��;"Gj�4!03 �O9�Fo7�� ��#�{��]'�<d�J���2�I����)�=���>Ey�cXL{\�B��B��}v =�_V-�>���]i􈸡x��u�"�5��[4�!l��v���eԌ��WXp� ��G�?�4�*m%C��G;>�+M�ݒ� �V[z�LkA�ô�*ל���m�����������d
���Q'[�cZ��Y�=�����/�������%�1j1�R���P����J�ߧ�d.=p�-�Z�����
yx��*��M�H_y8���6?�d�Rû�y���K������%Èig"��[��ҸE�	A���f@a�8����82���A�`2~ĥ~�
/jƴ�ϿM˘D&����*�d���Ej eT��8X�
ݲU%�:��f=K��Q�ͨ�{��Ŷڪ��i�r�a��;�p'ۿ
�ԲȺ�<�mH�v�|�՘(ѿ��dvn��B	+����Z���\�<^m��=�+�iB��Yri̲?���.�q;��Ȝ	��'�X���;D�;�ՀW�� ���qm�>��\Y/���\q��ťt;H��u��p=�ŗ��C�C�����~S�V���֡ t�Xʗ��Ԅ�.�	�<��h�����=|�B1��EuW��0�0��c��c��uSo�V�GbN�г$�M��7t�0��V��%	���zZ�ȇ[�m���sg��_�m����z��HV���:Bү@!}��8��^6X�ۮ>`)���W�Ä�+k'l���C�x#�)�RQ�ؗs9.�=��ڼ����(��1v�L�i�4�J���(�!m&�bQo��٠Ni[5��=��;5̆�|y��5{7�|�G)j���|!tn��K7�[<B�l�n0ʐN�g.�`~�~��g�Qm�c����nV��B	�G\m-lE|$LK���{���/�Z���R��h����7�j�⟮����4�.�cK��``N�ڈYRU蟎z�����������`L��YȲ�66�8���6�>��ŉ��ټ��B�6�a��2�Hl�RP�UMޥ�Vx�GʎWw٫�Cm ��B< _�;W�l��</3sŪ���`��E�n	�~����gd���16�r����1����Y�[-�C��Jո]�O��K��Tc�R_�d�d>#��UX� �)c4�fV������G
J��ŻK��A��r�1�/V \�����Nk#���<�s��K��d�pu؍bu	��&����?�`�d76�����4��A$~���H�>��q�'��r�c�3^ ���/Q�K��������Y8)�I�H���v�%��9�$R�V��y5����Ґ�*�!��i�:ﾗ���'�����!:�c�_���;���wB_��F�0D;��o����ԅ�;@�~�����V���A�B���ъ�T��o�. f�)��Z۠�V�5�`�U@��I���8����46�5�e�@�g(���I��P�����wr[Z�p��S�����J+ &�~�������r�xJ��VK
��e���u��Rhgϥ	OG*Y\A�ɱ�����8�噁Woڙ��kC%v:����&�?-4��B�+�@9K[����n���6�D�"[r@f_�}� �|�n�pW�4���:�q?mOy��L��ni�=ǉ����Դ	�!lՎ';$���/�I�H����
��*��j��3M���8,�"n��ǽ������ q�b���@M��_#�`��"M����,��"��c�����!���6��i�T3ъ��ѭ���X�O���S���m4q��b��g��L��.��.Q�5�7r�e9fh��{c�-����ݞ,x�I��~��E�Fh�,�#ͿNP�1*f�@���#�9�m�Uތ9Flk�Z
ʧ	��"^�τ����1#;��p�V/�ݝx��kkW�Jb�g3���Cίp�/��ӏ�k��F��'aNy�9P��^YL���ɣD웴����|qu�g�`�mQ�������+������������F.�w�S�v�u��rߢ�z�g,p$.iV��-|��VN�i��#pq$:�_;���+H��a%t��˵y߻I�[v���y�j�O���D[�H��P::�*�~��_U���ew�]%{�Yc�7E�?��%������$��R�r�	V7�YyF�����5�(���2�.44�a9072K�����\�ֹ+��;z�C���W0;yy	��bk�[�姞�j�o��,�R�x0���ow�P7
 ��%�AfndP���7�&��������{*=F�z��x�Ip�qS��GyBl����G�hJ-�lݜʽ�SO�	�D [���,�h��iȭ�?�Jx�9�|{�kqHjۢ��,�bf;��&ޚ�:�:=B�s�iʰJ�;%�vzG�	�Sh�g;��p��sr���B��f�g�4������5КH��ѼH ����:f�	���������26𵍗�*�/´��*O�zE-Uc	��;W�C`�?�!DHy�t���3�fS��a:@T��+I��E�����{�T�M�@m`ζ9���b���i��� !F:ǭz�0]ɷa��w(�}.tֱSO�g5��$��X�X�cF�X��w-�r^���µ��¼e;���P�����7����Эlu���A+�`�`�ƚpI~7���K���� �DV)zf`�z2�#u�h�<�5X�$��������&�$l�a�\вg^
^a�v�)�ږ�WX;G\U�7�K��2Uݴ���kW�-�{<�#� Ž�9����T��W�}�� �NH$��~���<2���z����wgQ�5衭lO?����mo2U63 ��@_3���!*����1��E�ޯ6������� ?]���%M��!r/L8fO#wo� $ϹU�.㊈{�#��A,�0�s�S�h�Ⱥ�����& �!���.�̆�3Ȥ�~�}�h���+<��i�~��G����I��§�l6����+b�_�' ���¢j.�"��#��u��>�$կ�<�Q�O/�CO��M�ZL��p��a�{� �M���Aj!��nh�B0��T�#���~
"s���&.���s�+m��Z��4�|����&��3��hNy�%P���hrA����:!~	I���A9p
�9VJ�1�B�~�떡7
�P��5*���m�WY���#�ء����u�O2푾O��Z>[x��r�q�O�u�04�M +Q��@�)��y���Z��]t��t�&���r�+J$z���:��'8����QmK8��\�Pg�n��ѐ�[JB�#�K�� �/x�1"���eEewd�~L��5+��pr�=�!I*K<���	����ISm�%~Y5$	��8h|�ۚƲ�U��$x���=ہn3s��1��W���=�^E���E
U��s�w��⇜���A�!X5\z�����h.�8q6tOE�tڡ����S{Q��r��*�ZS���Q뀉�|/�![�̅��w�/��4E�0�:�X�=>�Yn��=XM2b�wg���PZa2
Υ��PG4�Y٦���ƃt5��#Â&5�ע�þHh0��.��/w�͐�m���p�h�c��#V�w��܁$N�BiGr�w����� jY7�0"���Ǹ�7��Po7[>�y��|�7�����Y�΋��lc^F��i�rَ�p
4�Oߐ�]�GꭟWD\o�kj���>��A��� Pj[����z?�h�F���A�A0)��eD�C�2��S�3ʯ�w�XYO�y����'�To'&�����|�!Q7���V2�R魼֥��SN.� K�Ѿ%Ef��7�)P�[�,��p�q��cs�&����sNԽ/�Fr,;���m��⫷�?�C�x��/�`|���o3ռ_Y
����Rk�-�\�!no1	V�D�ε�
���HI�=Ҁ8~���-�,C��#p橓���`"��x�-t���:��83:X���}訙5�/3a1���7�H=Qs����y���+�Hn�B^62!�:�3�3�f�Zj@pl��bGmg���lK�e��2���Y���#���t�
i+w-z|W �&F�O���&��h><���>����!����W���<�h��U��Rd=5J�
�2�i,�_���xU�<w���E���R����<'w%�*PND�Lbi9�0�`Zؑ!���j�����J@�F3�wn�Bt�j�«�;��`�`צ&��[��y�W��.ڎ��^�?���Gr��
,��B��Ԛku�.*8����:;;к\��Jqj$���c�q'KΚ�����O]D/��C��
��q��ڎ������b��xU�B� /T���Fڡ��������\KH8?�m���E���ע�J�g����V@�<�D���2��a���F���/�iS��h��R~Oa�If�l����q�:f�4�$��P��l�P�I5��i�L�Y&CǨɳTfS k��v�{�)��th�p�V��>&k .���.Z��RMWD���[����)v�<;�rS��Xm�(�s�z0 �n�ML'�>��y�_��~��U�5���9�A�&sV�+
i씍[���(��;�����ߴ��^��F�h��q��[̅'n���� K�P_{V�<#��ݰ��TD`��	)�����&�}(��`]#?�Ұ����>�Dq	���,�⷇�a{Шqs���&��{�K���sg5πZ��8z*�����U���^U3k����a���U�A��YW�ؼ�����N����эb2w\u�W�N�ݼ��$} �������+��	���qF�*�oQSS0i��Qmp=��Y8 Q\��E5o7A�1L��{���;Y�|���'K�`�G���?�%��ZV(�DV�r���7�N��p]{����w.Ԋ(hZV���Tܥ�Ct��X���	�b�^��6q%:�i�x��vHu}�lWE ��} 

�&Z)�<`i�'A+��qNA��6��k��n�r �A��Y�/� a(�A�c����A��^���`�1�S��ۯ����"aG��{� :�"��N)OښI�@~~苴s�^鷲�?)N�\]����z�ºݺKpC;3(�Cq�OM.�q��kKhW�{�B��.�]����JB9�ĭf���B��.�����dV72}w�Ħ2jB�ܝ�O���Ǩ�X���$��Hh��w���
�S��=��![t�'�>f��V�4����b��+4�>s�I�����	,�?w-4�xRb�h8��'`�3�����b1{:���y���
6pb ��(����Z��6�u���tE�	��Ⱦ\�R3։x��*��j|�~"�?�2�@�pwy7S�=눿<b�>��i���x���a�U����&�V��7c����Zo������p+�t�uq2@��FM�yj1�״ם��qP,OU%PΡwK��^�u��Res�y*��q�+x�k��pD����*���z�c����a_zTcz<j�t�:ML]�w���(��|��LvL�:�Ngq�,���n�p�"a�FOz�=�&�$K�[�W巒nfʹ|G-����*0A� ��l����?`4��Ļ����nk��	�/��s�@=���G'�t������q����H�c��t0;L��M4���y��v�n{-̭<�NU`Q���ξ�5����q������ or�U�ff��x��>�b"w��;�yK�����ODX@A�AU$z{������*/V,~sȯ�L3�oh�F��R��2%�ǆ�:5_��EP�����UR�j�����@Ȍ/�����A�{�́,e�PD�)�u�(� �׎u&��i��[r�<�v���۽�p�%�8���a9�eQܷ�C�Eވ��FN���q]���ߙ�u���*�sVb�eZV|]IS.���{Q"�3'�����擱�g�!��������8��_}+�t$�,�%���C}���[Ƚ��)f�V&_JG~d�)�8�B�`(k��v��������wvX�L�Nji���,�w���dr��s��4��빴DXs� ��"Bt��B}rU��zN~fT�ٶ�g6*�8�^��bɰor[TH���*2�Y�r��/WX8�m{�o3����G������{F�[�pF2�R�ڲ�q�v,�$�S�=^���j�s��x�ɜ���)����j�O|TSR9����*SN�Ǒ�f9.FUrW�v[g?؞��L�f�/\��V�w�M.�e���3`��Z0�WNyMK\�4>��n!3��C0o��ܘӯ����"�e3��c�����$q�}w����^g<e ����R&��-��bFn��D�4W ����D�B�
�%:�4XO���T�������ځ��)��,�|�Ҫ���1g��пW�����p��Q����I�(���u[�ݷ�J�����x8շ���W9=7�Y�5�(�Qj���/g$)�[�@�UU���T�&wہ��dT\�<s��u�6U�}��,/�z���ͅV�0)�fe����&)⿲�]����B;7�\W�҃�)v�
E��n,
N�u�!�i����S��c��3)ʇ�.װ���ۣи�s��ns���#jH0��4�P��C
ü�0�Xt���y� ���)���v��9�zQ�*�U*�ʍ$�vn�	Ë\�9X��R|$�c+`X�3t{��^8$�=����O{S���p���4J�s���aUk���Q����0��� �_�.��	겢�PO�~�=����GՑv����	���+ާ!>�ɣ��$S8=F�3+!����9{��ʖ?��A���'�S"LM��#�/p`���4V��@���L2
p�	�Z�̸@�C�r�3���Ӱ�}��H��x���y*��ק��4�<�=eO@���A�A�J����A�������]GU�[$�=��=Kf?IB�:)��M ���H{�p���eуG'ɣ����{�IR5ե� v����	���Jd�+�G����VV��la�뎘�O�|T�����"7��:�B�7�|ht$�+�q��S8��`.�n^�FM�14
��h���κ��9�9��t�h���,�4�ck���E��"���Z��}aF�a����9�,uq `LYM*F=Aˤ��i�fE��%Dd�ĆMA�g`��7n������&��!�	2C �$��=A����J%A�]$��ý�
���|�U�}��կ-f�n��g�ks�9X�;��੍�C��m�C�F�Gy�'���:��QD�+�X�lu�=ōg�\G���E�i�LKv��!��п�o"�UY�䖍����9x����D��?��Are��n=��W@�V�i*Fٛ����X��2�?�%�-F�=Ú�i
�ɕZ�K3
#���N��fs��E�w��Zc���sK��_O=�^���7�[QJU��eq"؃UT�@��I%O3�@0r������|{�w�<"U�"����t3o�W�f���ٍ��<���5��M�ʚ2/�8�v�Oh���5[z�j+���Uk�\�G�*(��4S��@
:%�@�5�n���`�wN��A��P�iR�7��h���I,�p*�;�����H���Z!?t�
�D���f�*��֠LyQ�-"8���=5.�+~�\��yN�]*�y�*}�IfK>vT� v8� ���\}�A�g�.�|űj��u�	�ׯMJua�ff,�'v~ v�$�Tc���;�(�'�D�Q�����hJ푥I��
�x�\cc����� VI�'�$��~ ��O��ǐ �=Fj��;y����ܼGwv�	qa��	��V�<�s�CP� իZ�9Bs���x�rurKM��(�@�Q�o٩X����]��VN��/h�����+Mg�WWhyC�:Q�E�F9��Z�v��r����z�������� ���r�RMcՓfwV��8���-�'�l�a�E+f���/"�с�5��;e�I��T���K���>Ή�ñ����5���*�@�aڳv%�J5�I��q�6�d���5F�B��݈�9�W��~�u�Ώ���eX�/�+�ě\8u:�� Z�W�{�)����TΏi�6{��[E��7�h��3�x�YP���l��LN�ϼ�:����T:������8)>R���H!��c.���-��Y���'R��mň��ZҒ�4�SK�mm��b����%�ܽ�.��8��5`�f�-?�g����i�RQX���t�Q�#cϻ�M�>e�!���j؃�O
S}��^��U^:xç
�O��ɫ3�g(^ܥd���؉�v|̃�<�f��Aw$�K�8=s�q�䜫ҶD&��3�:��(�q+\����XL_�Ѧ6�"�9���#8�B}�»��+��t��v�0�1��$��f�s�e������!͝s��<� ��7>/x���� �@u�>Ri^�eEkKq|b͖�VL���O��CL<!Ԋ�QЎ�j�45J�J��X���vω����)/� �fSZR�m<]����w��� ���[a��!��܇�PD�N(_ ��d@����1�����ѯLK����4�=lx�<�Y��=,�x<N�O�5q���,G����zl��x�ob��.�|;R���?FH6Mx�6 �7�;�\w\����E��������K�ؔ�/��Iv��@5�*�a�y��kEĳPK�ԯ�B�Y�T�����*�Oݰ�)\Y�t�!��_	�0�7����{*�]�~"^z��]���2�k���u�sv��'wP��H)��I�u6F�O��������m�����'�����`�c���Jkƪ�q������\��L����]ɷ�(|"L�u��1�a�~�������ivW8DA���:�kw��?�/vv��q7\���}X���~���f�8/__u-�,|
]ɦ�``��l��e�Z���]^��g� ��Ю C�m�4=0�*?%�'�mH����r5J ���^VD�}+W�W}�V����;�Eiz��h�"E^��`�����8Pj�%\�\9�㐐`�nbuT4.o!�o�t,��(�f%�6v�K���%���+�����B�/�֮��߹��EGE���ڼ~ma\r����̠���j��^�>`s�\�l�<ߨ���`�3a=<���M��P��(@���`H������訓瓗�P;s������Lw������p���S�2��<+D�Ǜ�0����;xj[x�:��X� \�"D�t�����60z���~g�f�e�aOU�� .86v��|��Ifvv*�gYP�Ƭ����o_؁�5n���~'�H������T �~;b���>���X��W�u���:u4��Mq6,��ʒ(&��|�<�\�T����)�ٛU��I{ovy�}�J�W#�DDS�'�Vc��*8�J���h[AǒƧ��F�>���E5<���r?8�,u}�<��ȩ��w�������|C��������)7���W*�2��H&���F2%�e-=�j�TÎ)H��B�2����<N$1���G�u8KS,p�KHV�� I���MN'BY7b�<�q�3_ܻ��,�����[�p7�f��,:p��w��N��/bP-��n��~f_y�}~z���E�����$b�ؓq�X0a�p�!�'x
�$��0�Cn ˏ�?���������J&e��!h���/k�ʞк�ˊ54h�'h^�|�e,:�3Ʒ��z*���&��X�;��w�S2�k�`�0��I�R��G'��GK�{ͳ- M�>*{�ӿz��� ��([Pk�-8�0M���h+��e�H2����
2v�����Z���ȣ _|K~?���6���s���o��!Sw�Qߓ~4HH(2��%l�GY/oq~��|}ˎT���\,H��٭"30R���#=��Pi٬s��+��ڢ{��|>��V�ʇ�ɓV���"Z�/T��y�C �S����բN���@`N�f�o!ʸH�sd�Z;K��>2�jH�"p���|0)iG"���,�_��}�L#��ۧ���uI�i��d�i��5�T����G����q��U���OB���VY�-� ��m����f��P+�Oܹl�=�Q�e.�:��	s&�.��0�W,1�=�����=F���x�z�B��.�����w7v\�jjkQ��bSd�G���v[Kܮk�TY�)�tb.��]CN3%!��Їј·�`me繴�����Ȕg2z�fj}!����gQ?I����g��NԼD�Z`���ă2D혆�݂"�-�A^n�Q�v��w��Rj*��D�&/�eDL��?����E�%�ǓHp+7�7��_��O=D�;�p�
�{+�K��Ȫ�)�1��	������+�����m?�����(�ïw�ٯX����P����.��4=�E���m&h֢,�!0�:W�'�)�^�%�R5��Q�!j�ױ�O:��Y�G�_Y�ҏ$D��M;Sd�����E*��/�atl�5����V��ծ��V7�iw��ӫ�T`|��R��׮�ӑ���J/����}�����&N/B��5���9��;�`���z�{n��K��8� ��x�>_4 �!�h=
����-D��
b.�Q�M^ X�M>��m�ְ�uf��F���s8������Lo�6ڭLz�E����bC�"��5����d��� �'��@d s���
��n��͟��#��} �^l� �Z]�'��>·�������?w�a(	-_f�z�!?�"�p�t�'����\� IM۵ GI��0d�/����n=�r̽������>�	�� 4𢘽��G����m�lcm����7�EM��Ȟ�".ǫ?�Q����e���j(��Z�d��;�&�$�>u4J�T�����G*���1�6o��]@��N ��7�?�1�|���"���,�ڻ;;`�����JoPn?`�)@܋0�]Г7)M�bsUTu�/�*4�I�Q��C�܀c��$�[��dF�ǽ}�Kg��I��$�Ռ�X��u�-�)n5�д�i�5����])�=]��V���%�D�\DU�1�#_D㞰�TS6��;"�P�(R�~ QN�`-P�y��Ce���.�	�T���Ǧ�h�T|��t���ϞE��}�_�,�R��X����S%�O��&Ǚن��o�)�u2DnCx%�y�ٚ��4��8a��#���m�*Ey"��=�7�����[�]n=s�Ar��N��".�� ���Q)�pI��TABSQ�앐Ьn\A�*�C�e��1{��x�raQ��h������1yנ_?t@�7�A���py�v�/Ԅ<.e�e0/�,]e���Mg55��$t����U�m�<�K��ZI8ш��~r�'|�7��<�h��ê� j����o���eJqD�l^��B
u��Ғl�����m����m�Nd*�O���35�@��m*���%e~I�p�kO�)A)�s}��+F�;|��3��q��}(b����ښ���bJ�殻�&�	Rұ1�S�z��ϕ��.�)P�o���̣�K1F�8�0 ���	-�F����H���Z70]���i}; ��%jx`��Z�m?w/P��g��	�g�5b�%����ޛ|����k���n�6N��(�F���E���K+���įC�_�OƈIM��N��pn4�D�3!.$p�N8���:����.e�h����C���,�1`]E���%/	Q�G	_�9P<��gw�7�k�Ü������6�M���u�� �`a��� a\�΁�'2�t-XA�T,��>�4bQ�D��z�!b�U1�Sk7Y�I�KzFM*ŪـQ��&��c	������������$�����zJ�\�9nצ��FM�a�r���$��FhbL��_r�3���!�_&�AJl�8ܟ�}~N�Q ���AZ�N�@\4��]0�/��'�z��t,F�nIm�Q��)x�kK&�<4On�RM��Y�s˷���n��hZlS;_}��#�$5����c�7� /Xv�"C�Y�v$���gS���Y!���g���{�>k�[�%� ��t�O����X+A�տT��%�U���8���r"42�F�FĤG4� �?����紆Nh��D��;�sҤ�w����4P��I�x"�\��U�PeK̪��O��%�\3]�[.�q�슀�\Ã\�E��
y���s�1���2���75k/3V* e���m�� ����51�,��5䖂{�N�u��w�Nm$�O�N���u������i�~�f�uȫ$��8zŲ�d�����&x��䄷�1�m�����.����s�jJrb�4���-Ra�0ƁŞڕ#�z���笓�vTP�F&gܤf<�f>����ҍiDu�G��q+du�$���/������� Sf���t7�mĈ������9,biӣ�_��U�*��//����� �"&F�k��I�z�� �l���"B22pއ���!4�
�.��f��a�`�E¦3,f	-M�s�P�:ipDὼބ����O���<��F��(p���rӫm�c����AIQ�B�=�4����Ź%�v$9�l/�%?�|#���'�٢J^ p��m跗�1c/�ȡ�1Y����\��>���s��0�@�j��]��%t�npW��d��B�1y�f127�<�آc�N�];.\5�l��aN����X&�Gr��J/�~���t+��
��:ic�UF�hg��ȱ����MTu�^q�� �*՟L$�(�uy��h��4���7�����̐�/N,!3�Tɩ�_U#��r���UA��4����PN�ju�����}������Q'��P��q 
�W��\*�	Ku�K������&����.����}��*΄#�H�JNg��P`Lc�-����5o�`��l���m5Y����T�4�̛3j5��r���`Sl�h���̽�D�����LM�^n�st	:K�Ƨj%"�r�#��ܖ�c3�J#$�HQӛ��Y�Grecg̍{v��0��j?O�G����q�t���71�CR�!Lb�0}�C�^�XS��h���dz�iU2�?.M�n7A}Swh��$T��C%�l��ʦ�OH�+�YE�U�k���B<[B�8��c�ch�8�A��{+��#���(I�~Ԁ�L鶛�KIZ��[��I9k�} ��U�-���Iģ� �P�ݕ������1{@�}M �Y���/ѹv��.�1�J�!~�j"f�g��ڈ04ϚK��+x�R�ʛLU��|F¦�.-���}㩜�2<6/�Ui�������"-�fȽa�"j2mO�ne2�69���r��UҤ߳N麂�! fП&�ӌ��C04#�\���I��f)!y�s���Y"�� �2��AO37����x�C�\˯e�����g��ZFZR,7�򑕔R��ꚴ�y�p�6TLI;�M3�I���I��ZX$�Y\L��0�{�#�����W~<-	4��H�q�/�V+�:��X=�	����ۼ�}��76W_�c�bͰw�o ��gmȥ��2Kl�K8�=,���X}���v��e<ٗ�*�g�NĂ��t�3O��#>
7�9��b�@��M���]+�1���!b�k:�OP���U��(���IجJ�/B���׈x7u(),�r����J{�
6�s��Rb�+�^�ҷ�Z	6��Ϸ��Z&ڛdC�
q�
��U��A��˯���3�C��a;T�v����U�ƅ�LeO]�,��*�4��n�b�җ���Hn���:�X3����F�l�܁�{Cx��c^[��d���QA�~&��j��#4��9���̆Tg���v�V�W�)���V�g��^-i��I��]�5�-g�y̛���ĢX<�dLNJ4��7�nU)�'�<�M��Y( �^����#��s�3ٔ�N�Z06��xBp����qt�z��'3
i�֬i�*�z����$-�Q�?���0��T��=��^4�0C�.LƉ��8�����+�D��D����k���u�ܢ6��C#�R��!ZB!���vN$�$��$��.x(j�����0�V�sk=� ��y+��4�@H�
I2��L��}�e*�a�U�'p)�F�����n靘@��*��i�N��$�p|t ���6m��Jx7q�y�fMdЏ}x����/vq�1]����Em��ёR�O�zJC\d-s֡�Fӧ�����x���P_	���С&�cE��5h�BmJ�1��)��7���r7򪷶�o�BK���{W]J.�I;�CacS�/�ڷ&�&y�ܺ�y'��{S[����x��D�sO4Rk��E}�����8t�>����e#�廒tǨ49S�3��>M�������:�Z(�]���XL;g�@��q�R����R$��I���}�:��X�u����[FWoX$e�f��u��觳Z��bA��/{�\-Ը��Zyȇ�J����?�.\s�@,�V�0��F��b��`4���e���s=������=��/A��g�gو7R����� ��,l@�We.�L�4�Q��IO[�w�Q46�1� 㣜5q�ǹ:K������ ����$�/�����g��ۓ�*�p;jE���ն�3!�����׊�ᮔ�Y|?�~�gUX���;8/��(���B	�%�&�fZO��b.4��Z$S���N[~5RI���|�w����=�.1F�陵B�%��s^I7�t��2l;��	�j�9<�S	��b��ܼ�u�-=����S��Z����ج���UEch���7Ɲ����I��������uҚ����?f`u�bU�4-|�-��}��ڄ�៴���fQ���&���X���N��M��I�ɟק�)�����h��Z�\� �6����e�!e0��Nӂ,���	h6+2�`7�ω��q� Gj�eW�y]�l���ޛ��YRю�h��1�����c�)|Q��	��/�vڡ����C�a����ez��Z�z����p�Ib%�4�n.t\�v��3� �e]�LխW�@���q�N�I��E�)3�o�ϒ�N��y�zGE�f�(k��+}�<�c�db�HD�z�_��l��҉'�ޅ k���>�B�2^N�'�B�@m5�tzz��`�Z,k�/�������X���Qr#{�����*r����,���B�[FDԃ��.H���]޸�6<���M�5I�����1ƨ�_���d��v6l�.��'�<=f��:I��G�b�vK`��7�JX4�Iy�(�`��΃��I�snt/����,�[���<�yD��������yQˑ���Z'_%�/�@���F��M��v�m$�����4��[�� �9wW ~�I^�P����ֽ]݌��B��_/9gN��ơ'h�̙L<��Xw�ֲ��%[O6�J�^r���*xh�~�ʄ)~c��	o�U'�,���r"ƢU>�s��k�}����J6x����S�[�h�S��w�E8�V)�$�]#�TڌF�+}]�����=R0�/��D8ĄY�H����ҫ��|������dY[��0��g$s���I^�iHL�8د+80i�A0��>݃˕%4�X�$�r�Zm ��v2�����	O���77��>��WG�;\�.e�!���*��|t�7�DD/��@��6q9�}ɓ�p�ʥ�W��ܐa7����?h؀q�oxǈ��Xl4�H��j�m!}����+�">�s��]��10��-���x=}����� ^�ݺv�U{4����u��[h.�%��$e	:�R�mE�Co\G�����M������e*Q��ǭ���Z���y!��a:�̏�,�\h�������q�.�}P>�(F�4��`f����i�As(��ڜ�]�7�����$�̼�� ���0`͡?�^ߛ�M(�t�CEhF�Z�{����7��� f��A�� ��X�R�h����OS1�#D�>F��/�.0]<�"p��8�o��6�Zі4������*�<� ڊ��n�]q�<�Mw�O\35�]�D�n*�6!]]5�,#���{� �$�|�;^�
��"r�C�������8��W�ړ���q�q��ּgo�YR��7|L�6�q�9����d��;�&����@�� �頺ʤ���l��|��!���?h�;V�}G�H���J�g��7����_�C�='�����5R��v��*��W�g��>��UY�gV�� ].;��`��M3��g�&�]}�`�9Ɛ����O@�ʌ�M<c�&^�
:�*M) ]\�\%�=e�����:�uj����}UY���a���s|+#�X?�[�A����(۔$e���B��� ��X�o��7��h��A�Cf��G;J>��;�ő�|��b2AG���:�N}�����~.�Ula�m�=�ɓ�V�{�D ��U6�6�xy_��<^z*t6p�oUC���kuE�pƘ����->�
�;�s�0,��ڹ�9���8������R��B����U�Hq�� �o>6	���
���c�p@Y�E���*��}����6
�+ժ��1C�q["�0�s�W��*�^S�Ɔ��I���g�Fy�.ப�g�%���Kx�R�R��OOg0%9�g��٫� ���aT��?}�1z�J�*����?x��t��E��q?�
}�1�7�ͩ�Q;fu*���o�2� �_�G���Uky�,ƥ���0*�l��Fv@�W�~�*�^_�h,���ig��j��$F�n�$�W������#�Y�q��I�Hӂ��Ͱ+L(�Y#2���2�����*|}6�%���<p�͑�C ",�G���n��ZT����Ὓ˗_t�)"><C!W�����tC�F��h0����H��q]�g�%vg�|$�Z�P7S����ʱ��`���Q&�;h�������]�^�1����}����Mn��#�Y��CW�.��������B�iG��,\�ﵩ��#��8ڂ�V75���Nm��>S�8�4�i�؟V1��T9���R�'X��⢭�_|��f��q�%������&@Q??I+1JC�\N�q���}���*wW&�Z��Sˍm�n�z@�H���ɬ�pS��	ډ�%��8P;��s�d�*$͍D��Tݵ��&�̱C191���5:�Y�� �V�"=�NQ�>_w�Q���b�1{.�p	ּ xR�Tۦ3�0�gz�DB�n�?]������l~xD�JE{�V�����hH]M���e��dhY��: ���h'��{�	���H����̚0¹�Ō��PC�M�0�ņ����S�:�9u�|����D��Mw����zi�A �q�����@M��d�)|oƜ���h�`A[�a�Y�S8Uz�rZ�:)����#�T��}��o�ݽ/;e��� Y@B�$BnG�j��@!yE=���>�V�X/	7sˍ>p�gU(�զ�r�5�BS�*y$�*#a��AJ�-��m�4OE<�Lt�mW
A��3���+�No�-fH) ��I� �_�h�B(؊��Z�Q1��3�%�3(�������1��i��E�hs�U�~Y;󉛲*T�<��~��F$�4K����`�I:)�j{;da[{�~������ș���k�>���t��c-��>�&������e��ń�:��#Ҩ�~�q5��� �L����(�p{0Ka�n��P��)����������8�I��D�MI��)a�h!��=�ni��v4蟕��}���[�֕��,������;�H����:n���e���sLL�g�(�2��yۻ�#X��,	9�sj}�!���춋1��s?D[ܵ����Hp+:c�	��"����ٕ����Okj�nD������Lal�Z�<���#Ck��8�b���Pv�IG1��6Ś�
�(�<e�{m�C��J;���U(Zu�+�3�ϝ���Ԥ���a���Y��*-������!��HI
�f닫$;KWˀ����#\�4Ҡ���o�8��h��q��k�c��<����)��2����*U�H'
���d�Q¡ I�y�b�!͆��]�#����𻽾�M��d���l=Q,(΅��ë�2vŭ��%2%���BbO��̙,�B��3&9���CGƉ��N�o�l�6������f��~xכib�ɻL�,��'�v�P" �dy�S��K\�.�Mz]�w+��U`�-~��STD��%ft��3��R����q��CP�:p��� G[�VO�$��k媡�ѿ�vd�ƒ�Z�	�^��$��z.�X��O�Ԅz?�M�
l�������<~\�]�����V�
z]�BIlPs�n��Ɋ�'�[;K�U��9Ƙ���uj�Y"��A�� .Ű��X���JSu��*E���m���w�[���bZ1r���rݍ���kbNw+xc*��*f�K�Ne;mwo��/[`�����ı���Yd�����k�o���������}�4��7JY�4�s��{6�}BFIf��Q����ܴ�~�$�����)�ڒ,�p�A��]a׏�ve�lV�̐�v#>��A�pD1_ǘ�����H�?��k��]3	$��T@�Κ�Ε��X���.
y�:Fx�-v�̢��Įw=�����|� �o������{��f��B���}����g����:�a�=�I�%��`����Nb���C5���aJ����+���L$R�e�Oqm�7҇�����f7l+�,	�W���������g@F�=^e�g�L�ɡ��@U�a�doz��7!������+<�2�O�S�E`�-�]|Q�fe�y�f- ��.�u ���W����h�1�b�9)��"s �j��/�}���2����:��𜪼k�]،v�@6��M��=oK袲F0�.n�U�HI��R�z��}���:��%��q	�sNro���|��m�m��-��\m�Vt����
%��(��v��M_���~<�b����H�vkT����Gl�����9ok�]N�nw2��ҟ����v�\�4G���\*�Y{jc�#�Z{�_�P�E��U+kN@f�XO�����l�Pdi�^�����r���*�}��^>�f�)�P�!�D'��7�4���$�^7=A9�R���1k�d���dI�_k�[
w�q�6��T��{���Ry3��P�\҇�%�5O�xl�ħ2n�J���U��U>�I�Q��`��>6�I5���\��91��W�F���pӡ	�T���^��ӄd���`�%Ј�� �_) R�̷�����닦�4\T��M��/ѕO����{ր,���X����!��3�z� N*>^����u-�a��N�������6`���~�P��f����B6�D٩�A�]��p���yXڋ�`�\r���5�2$ݚ�__ՑY��D� o~�X;wI|tx0��;FҭB������ ~����Ҧ\¸���i�m)@����m~}f�v�GU��	�L����*)���4�"AL�M��31���~5��G�ud0L����-���E��B���F1�g����A�~v56�v{���##���fRkI���u.i����[����:
zPx���,ǽ�Xwt��q����^pyV65/q�}1�^��c�����el���J�����cY��v�=8�Y��)��������WZM��#;�Z�j�I��9w8hpg���(d?a�s%��ʪ<����{��\EREj6�e�%���(y�g������B�*�Gr��RU��l;�	�c���\͵w�g��n��U���M��,��b��Z@j�`�<�t<��VQ�p�j����������T��w�@&,\~ %�i^�g,����(�찏^�2ߧ&������U=�:?4~-�p�Ұ����=���%0�B��?�w@�c�B��c.�/�]B��8zӠ�䦼I��Q�?��B)"#gI��-�<��m$e�q i�@�m�7�.
�=b�w���v�����^���QUɲݗd�BK��d*��n�7���<y�)&�P��X��ǯ���cϼė ��Ѿ��JPkY�<d�w�a-pS�O	��|""`�?M-!���|�UFp^-���ө� >�Cs+z-��)1=`-������WOߦݲN��U��@uyD|Hju;rI���@�YV�E�[W\IǥE�"�
}��[-��U����E�*��|0x
|�/�q���Sw�h]�ǩ�N���w�����OP���@P�f�_}_����g���[�ne�.:�6�[4�L!\]ʪ�}�'F�&�c�%WÅ���s�z�,��}
U���qcZ6o��S���EÑ^���r�'���#cư�)�3�c����r^����_Q�h:�f�<���{��n�ٜ'DFX�7�=�1;
�%B%a2��0�ԏ/\�$�`g7��� N2z`�<+��w�,���s[��&���\���o��H��F����%$v�e��j	N>`��!�_]>�qR��i_������K�9���n�:�S�w�F�&�������o�K���<{��l�]o�ڍ�]��v��<s�	~To��� ^ph#�'IE�I#��_��-���A�#g�5¨��U�E�u*�6���q~)u�Y3V-R�	G!�zX�iG[�兦���_�Կ�U��H�[�7D��"0���~��4d�N]zH�f�5�ь��
MtD8��~N�PN��]Y����2 Z�������j���$�u���Sk!���� �^w�9"J�?�,��WM{����*z6"/"�����("�:FTD��(ʧ����N��:c���`��$�b�)6]^(hO�j��g��U^��g%�@"��2�e�q�Bg{���4�N�urƢcc����r�+g��⍛9�w�C�	{6��6��묃���z������3��2��g�r�L{:�����\�e�ݤ������1�eQJ4&[���Lw���s�i�ޭxy�/m$�'MSӚ?Ξb=l�H{�q�
Z����o%�;Z$� �PK�� 碂�Y̀��$ǉ�u9(3��O����?��!�AhpC�
W3�s=/�nl��?sx���ׁA�C��$wZ�C��@!�|O"˵u7�E�DLï��+DuJ4�K�by�
Ejs�������QdNQ.����j�����?9��LjlU��	'�, ��y�j^mg�4�:;�I��fT2��@����#;�_��-$*S�y}u��\�݉�gJ=�	q<b�w ��i�D��
��z�s8e�|�k�ʐs����μ"�Ȯ�L�1Tж�%6�x����4�`�V��!
3��������h��3z��_��^�
hG��+�cO¶��$i���ؖ�)���R���>�Ž|��Y+%l�̍�&��������A���0�+-�(X�*l�c�pC�O��v3��E����S"�	��S�^�C�?$�`{<����f��;^�46�U`�`�
�-&��}������ӏ�n�i������Pd�S���"�����2(?��9*{��J¸�ڝC)���j�k�UJ���ttL��XKY  W����6��3�`_�8Zpv�w^�O����s�8Z9�6�k!ؙ:;��Ù� y<q���XQ!W�i�5@uR�x�c�l��X���k�s&��zg�O
�
�$�,�����,$��ԫW���b�I��FMU��Z��$�]���"J�2=�[�����8ٴA�k�g�'����ر�n��d�K�r&v�h�Сr�
�R˘�����Bޓ�$8v�,�8�O Uگ�m> �@~�-�K�g8YEy�Ӣ��ŝJ�66��e��!�ZWV��7$��w/0]�`1K�P�	�&�У@5��#O�;��+���O0_Y�J���koV��o�.ͧX�\�[���i��S�Kv��CaXq<���{��G�*�`�oJ�9
�d���6�l����J�S^i�ۘ=j�&<�2j�>�� G�J�\����cL��Wo uq��/9�hO�4d�V1n�C������ܺ4i*ƣm=7k#dq��da�&}��E�%8�,L�|!k�L"�����,�3���N}���e�����< �ԡ)8EP\�֊�$��dT���S���R�ca�N�'�1�D�A~A��E!�T1G5�O>>�u p�L�)�g����#��#׽l��\�zTuGU�j��*�	8�A(x֢ހ����B�1=R�`�a��ȉQ�wwD��.� $l�Ϗ?tݴ��G�=
�,�&.��Fܐ\~�J�����G(�K�٧q�L�y�ro�,?.�?������7Z⺖Yf�{��,�6}lK���J�@wI��i��#]+�m���O%�Av��t˒9Y�Q���FfW��䕥�u��["T8�k�1��|@�L�R�F5T�a9�('l��WĜW�jt*����l�ݎW7���EWP��c{�0�p���v��d�p��!��]���'��
$���d|�PٗMxT+]檞i*H�!U��ܞ���X���|Z(.x�k"Y�(��m�X�����Z!��I�uD��$突6�-&���+9��� pp��wA(��8�g8�.W�oH�Y��W�3qgT�so�&ǽy7u��|ѽ����Y2����??���>�%��z��)���ک���Ή0��OT@�)y��@�kwb,##[��TxUؒ��_�%�V�bꖸ��n�t /&�C��T��r����(͛���2K�e1Oq� Re1�wݞ�X�)w��nȟs�&&����hzd���>�Y��f-�����Viȣ��w;�r.�� ~yxU�Y+�[1��O���[v�|hYe��$ 1Y�����2U/�	uC@h��H��i����6j��P$��\u��{�g���(^�>�#��?Σy�=�O]�;��U�N�b����/Lg�E�}z��a�T��J��Y�P_/��e���{y��zqe!�	z����B뱎T�GU|���7�7l\�v�ꔄHlؐ4�_�u^?�"���h��:�͋�J�-��m�.������`
��9�@Ȳs 5{�Q�nCB�ZA�'�k.���0r9��r�����&�j��m�2lW��H�)f	�N[�L��Gx�4ŝ`![=5�h� �o�j�����s��J��a�n2d�,�}�fg�?o�L0FiP�hA���#z�[���Q��!@%�B���b�jE��)'�^S��af�f���X1]6a�3���/�͜l���f���xtL���
lLm;m��N���ނMp�r>>��J�k���,&~xw@��'Ͽ+{�<M���� kH^T_���ҫ��X�fC�7ʁ��h� ��.E��	��-�T�4�?	� �K`��st�=Y0)�m� �aUKg�����4w�u���[����1�� >��-*rK��\��vɫi���~���O�ܸ�9�l����azC���0��ZP�{͂��^�a!� 5�,d4�K���R$y+G�6U9�d�\&3��sW�_�޴�O��K3+���ZKX�]��,
�ZG~�>�LjU�0�N}���~e�U�Ҁ�U�&S��*�� 9�������,K�+jh�L֤hB�����"��������᤯$�"��R��J?dR��ec0�V����iu�ܼ��U�p>��l�9+�l�T*�8��}M���qO���a��9B꘳�A��Lϼ�g���Ƙ���9G2"j�H��9�6k�I$�eZ��W6(�+?�J������Zs�B`Bv����~���_I�9�%W 2&�ٙu�w"��.K19���r�(��Idf��0��<b𳆑nJ�G�i|4C�ܿ_2��*gCÜ�2+�
5�=kp��K�0�-mL�I՝��~=�d-uv���N��Nv��@}�O,�5%}5!��YR��9�&��bcg������j�IN
��8����a�Ob��Šc��ϫbr�IB@*Q��5���1̅�4�R�fYd�8�k�*)5�$bƜ���N������B���-�b�t2r�`O\�>&�<�z��=R�]��|U�<�[؝��>{�B�n;��y>�8mcZs��Μ)��J�$ρ�P��b�)3�;��L^�z��}cu���P(��^�$�s�Xȴ��Y;�<vp��d�2�0��t+��a�@O�ד;��N�ȹ�%�J:�g� s��+&��?0�C�_
�j����9��"~j�uь�z��%g"%*�SqWK���tZ���<��i���w����J�����ƺRCF��s�p�� _Mi�8iP(����6=�ht~���B�T�ʼ�:��0�RP��j�\[svW5�\{�y_ �_�O��~�M�%jS)�����	ͰXگ[fL��"<@�1��jY�&�>����Ag����?�/d��4�~����/`�퇁j�<F�U �������0�"�}6g�=X/wB��GM�8�|~���؊�`�������7�Ž����ϑ�[QZ�׊�7Ni�t��c�=�<���������0'���@iVK�:�ǋ��(y�y'a?���,��`�e����d:�t���:����u����ͨ���Ayb=tp��9E5|i���Hc(�}�󞏢�/3�!^7A#��*�"8�z�!k:��^p����x��I@Ӓi��4�G���y��o]V��,���ws�jf�=j}eo��@?΃�������ճ8�qr�_S~}���
�l?T=	c��P�R�]k2��"�cٟ���J���Z�)h<�V�l�"zb��HJ���&�L<�d<�[��A̹�PӚ�3q�JXd�U&X�K���a�������P�I,�GA��!���9�j˷g͓�M����r�Q��*��a���u��|-@�2�A�u�Y��kn軐��LB",h7,�S;x�T7��ڵ1�4��X��|-A�����u*��k���^Bv�e�"�h�uc�	��:���t��]����̀���80Z��8����.O>�&G�׻ьu/Te{Y��z��#*h{�� 8�c�7��������V���+ڟ��|�2&P���F��%�fu�{�U���V����A��R;�h�V�2M9�o�_��&'6e����b��z'a��  HbVs��)a���y�`��q���U�?����>sJ�+7�=}�P	5��H9pa)gV����]�c��*ǿ��ز���3��Y�y��G�9�<�t��eW��_��Y
A,3�\}�h��j<�U�����cO4ڔg+$���' ���༰Y����#�'�%I/$,E�-[`���B�H�:��x�ٳOZ[&iX�|>�8�n�ڤ���p)�%S��ܿ���X��n���e/������SJ��t�.��Vޚή���^!�O�kp��(b��g���J�v]�#u��^�gv�bz��_�/��m�c��6ZЏ�l��20n5���\б�+P�%��
�P'Ob�<H:�`.)f-/���e��]���Sfz���[�w�/���p'�+�u�Q?5�(�o/���������V�e��O9���|��ȁ��&γJ]T��W���"��w�R@��F����%,�x��*/Jң����p�_�D� �O���@h*��d�v��
a����-_\r�HP>����C����0��fU�`u�A�<]E��XE�^��B���a����}�����0�0Zj��#��r�J�@��;~#1A��DP/�~���$TV�-���:����] �@S��}�U��}�U��������\/�%�o�X�U��:���0�\m�ŵ�;&bxYШ<��QG�SyI�CD�xy�/��LCQ�d�lܪ����!0;>k�;ƕ�˯x�#�'��\���*j�b^a�u�i����9�C�}e����5с��5�ݒ�dB)��Ѫ�6�"��V�-ʿi=������I��t7�K;q����I���1�:���e<?h5rom������c������K�p������@��+�Ⱥ.��c�e(�E�����h�p�������m^Ml�ǂ����R��`�}�o�1n�6GQ�o;})
����/�Y�g���~�/dٯ���$s���}%��v7�}8���Ak�x��L��3auS�䘆1 �b�P��_�:&���;Djht�j�C_�q�LFͬP��tlS��BG�I�i���X����S1�V>���zmo��
�GNַJ�Y�����}����pʲ��"-�������wA����q���\����ynҟ;#��\�z����RՊ���V�	[��w��,޵��× ���o?�I}b��q�j��_	�óȸ����!>I)U~��τ�~���cx�gw�:i�n2~��u���Y49b���dq�,��U&zOt`E��x�Ϟz*Vh��.`h���G�$�{_\Gݓ BAT!��J�+<��Y���4����/_%"c'����կm6<[��R���gq�'�$��Kj2`q����C�gUX;<�q�r�Bf�v/�}�b7�<���� �;]�#"c�����}��e�	� �Md�oL���^4�A?Y�ޙG�8���l�d��|�9n\��.z���V��7Ka��&O��᫤4l�Ar?���m���l�lD	e�'�a�$֌A���P{S!Q������3P�
چ�ڊTp��}�"�������MCs&Q����|=Gͳ��lř+_��ٰ����r1��9�v�O�%���� ����?~`g�
�� ,mfI?��ts84����
����_����HI0%��ܴ�� \�*�a�ь7�/�ӄ��#Ŗ��K-�9�y��.��Y�|yN-��Z��$P6diá���(�����:h�B�<&&�d�n7� `	���Z��:#���� �UvBо��>ro[���H��#��h�^� JL* n��14�7G �ך�M�a��n
�����
YA�enO$�0O˅\�8��K1G7$�"S( ����{�� �A�L|����׺����r�����"����V���}@���{(0��XA�NK�� �`�pyO��d#D�C?��VR(NVz
+��Ҏ����z�t8��2�g��d��@��^A���H��r�}޾+��1���Cc�O��3Q�og�C.�mwZ[���HG������Ѽ.�&���&)(��ɻ�e�y�FXG�㴋mw�1�6=��_ޯ��,�[�����9L��F䠗��
h�מ��D�岮�h�J�R��#��I�BvJf�ugR���c���B�W,q����C+b!v/�
l������Qڬ+���!��Kw�wRQL�[��r��w͹Ķ�T�N&�w���Ql�]�>ه٧BV^HQ�r7�\�w���{�kD�o?�;��,�}?(��mq}�1 H� ���B[j6�epʑ#b_��}	�H
��ƙ�=����<KV�k���Lry��m�V[nш�ɢx>�"���JW��BZě��䈀��N<U����gO�I��_�-Q\=��}gB8���t�|Mb�ǹ�6��O+QH�(&f:i��pT_�՚��Ʋ��Mln.r0@u�����a�h�R�ͳ��2�"(�U�~�v�s�D�/2)��7�-9�{��������;�'#�o��c��q\F"V��,��y����H3�~+�{=>\Ĺ�����5�A�����R�?(b��Ԟ�k�M�s���%��|��4X{|� _
F�7�Cl���+��D�Q��Ňu�D�����aA	�Yi�M����=+�fd��e��b��gT'\�zhSK����[b�C(E�Ú�'�KT��Y��D������(�f��ԣ��]��@��ifk鮈���@tl�S�����g�)�ѵ��->|i��ȣ@��P�����:�z�����t����\l��iv�u���`�B�lH�?
��s_�>�R�J��f��_I�e�xQ����-�~a���I�xi@d#�m~����<�|��Ӥ���⩄󱬃�qD����8U�jp#P�ğY�3�X��{���|�h����G���8��*�dGl� ?��<s�0�h��<8���,���ʖ�cd�-�=��M%;9n\�v�{0��񃝕7�q>�����#�J��yu�,��E�TV��䱙\�%(�����*�ƴ]ᱤ�4�aD�|%�U3H8��:Cܯ�r#�Dt���pWe�V�11O����5$�������.���朌�[��F��1��>����i;�R|�ɻ��UF��>X�TGX;���v��A������G�n �e�}����NT�/7��f:r]	V#(�����dq��Ħʝȫ���{�Wy)�N��v��@���{l[Gͨ6y���/ۄ�:xD��� ����v�V�
�X���*8#�G���0^%%��Q|&R?�&����3���'�U���h{֎��7z_*lY6;!�M�c_jdg��K�
>�1|֝)��f�y���Q�$Y3�� 2rJi�l����4��<����]{��8ma��*�:)|��u��O�&?�c�}4Dq���'�e�����!��9��G�j����y���4�f?ar�K��C�Y�HFߓ�5@��%ܢ�`BתO�.2�J����z�V�3�뙎|Őz��g��뀤�b����C�ϓC�2W�8�*>�#����ۜ,�f"~#�DI�h}�Q�|�[���.�M�$P������F�N�@�ʹ���mG���^�5�ZY� Q,��]X��M=s.Q�P���z��Eߧ07�r8B��(aq�F�_��pBoVa(X:�����R�w�9 ��f74=}��5�,;=UKd�j:$�Y~�*+sIK��З�����<̅w��?��ӷ�C��,,	���"��9E]��&@�P��CF��m"�zM�J�ڽN��U���޼�q���L.�Xyc�����/>I��z\&*Wj�v{`�#uI�̀KԢ�6����ڌ��Z�
셆�FE�ie��TI��ńz�>(֜�yEa����UR�	?Ǆ�W./ܑg$��/�hX�0�8]L��������Ȱ�ٗ��%L�}���pCN���-m@��:}�{�k0�Fb����$���v�ΥprP��:5��i�&Z�˫d�cc�=�8�䦸�����YĘ�7��Fp�Y�
�r"%	�P8AS��2���
�z����{G��z����4	��?�JQ���J�]cӍO�56[��7������
�U�C���Z��fU�&��?1�����mm��S9�k�a`ۚ�)�4��m���T�u��ׇ�,�
N(�����i-�	`�Rn�N�+ 1����3��
w2
�3�X���1��0���{Hd�c�PZ��'=���ݘ:����0Rۂ�l�ݚ���q�s��;Wm� S�]�ez3�13S���
2�oj��~���XG��+<c���I���6��p��E.�.%����,��`����i}`�Dp#$���L��sM�x��+`
�Q��:BK H��t$W���Ňx=8�
���}��W�A���#��tp]�C�7�d�W��H��ԗe�j
��)��ٖC�[�������������ai��Y����Dsg(z+mfUP"|̩��xR6���A{�Eg>c*�\|fC
r^�7���X&zk	��t�g�)��y�?4� �6�UJ����z���y�H�	oK3�a&�L���~5��0���(h�����	g��-�T���K�uul|�Aڮ��n�Q� (i;<v!<�3��N b��o"7�X��`�P�0�9qh��Y��>�tƣ9�n9��]G�j����ˤ�IX���PUf�X�添iI��F"& ��Y S$O���[@N/3x!B���2��P�>4(,����'io�}�z9_�ˮ�̝�� ��p�c��K\��nQ���:�2��kې!g/�7�a��:|k��V�Ք�,Y���!rmN�.ѧՑU7
-�Xc>3��֎��-c�(�@k�(��5�����=h�:��V�֤��k׾p�����ĸ��XD��Me0f�6[�&6�zԷ�vI�� %�[n�Ep�rν��|9��_+�,��1�j���ɲN��,N�?�.��[�~�1)���s�S�s7��Y=[�<�F��;_�ևA��.������&��J�����`}b"u����4�Q5�_�p�h�2fk��\����z}�=ʶτ�g^6=���G!�P�R튵5?��+�4J"�r�;Hī�W�L������3�f��W��8x�r��Q�0��J>H�?�����g:j}�pD��f1O��kׅȠW@@�/)D���(�W�DC���c#��'S�����U1M ��R�B�O�ֲy�9#�}�n@�N��6�zVw����~�jt#T�o╦�
Rp���"S{�NyA+rfǣm4�s3�:�[G7��?j�
6cL�ɢ�"���]���gxU$����zC����`O-�T�&�&�sS�v�u,��Ֆ����B���̯#�Ō�n�*8�9϶��3����pQ\)
7�}��������L(�-l������<`��#~vs[ԍ:|�r=���z������|�g'�����R}R��бa]A�Fb�rX�|ʑ	C�&�� �'��|!�%�I`��E����/�K=�y���6s^_Ʃ�����!��L�-����޽.M7x�K�4�ҿ>��N�n�&�I6�f���H2���ָ��R�@!USܶ��ZE\C]Kuox�Q�� ye��mn�u=��9p�i�i��{�=������V�����`픨9�H@QlD6ʠ�~�N
���/�`OX\��ٗ�ݶM���7�5��.|o�A����	?
�]Z�"�Q�'A�3�>�؛�7^; B�ԯY��ӷ���H�R�������d1"�j�"On�c�f�!t00*"�S�@�!���d"�;g�xObBaH��$3��� �����`��vT�I"?$��qI��	Ɇ������|��I�מn�+la;f3��NPԥ�ƙp4�H����)`(XS)���tݍ'�./�c�=	��<�"<�*���BWU^��V Э� .����$�D;�	ޜr,��J�;��0��c^�]μ���IsߎņWt��٣"�5���+���sR;���f<�z²=��ޣP�%L�*�,���"U��F��R���������c䫙Jwwz�dmIG�Ia�U�z�vڒ�!T�C�����~���Oq.��{�XeĄ��Ǻ�[P56����oR�Xj�X���M��ٓ��p��b��n��������x�W�j��7)R��i����6|�t�toP���& >H$[��۲k���2��n�o*��a��oBC�:��Q�(��_�����,>���M]���*&�%`ݠ��������=OQ��A%T|pڎ����dJ����y�Ɨ�W9��S�F���L�o��T�5t�6 >�4q=r�E���|�;�:
hr���۟���6;�x�F:tS���j��܌M�g"�j@��}�6��P`b�mf��4��.�Fl|�G�r���R;w���մ֦Y>_,EE
&����u�k��$V�s�ư�s��Ϡ������$C��QL��Z� ��co�m�u5�Sq�	�&�ߐ�B�����]K��?���7���yn8�}�(��H�4�(����K|��l ���3[��}��$b��/@2>���.t�G�����e���T��s�D��cځJ��T��_��r�JmM�:�a�⧓mj���<
�hz��D��E�n���ğXt@/5��_��|c����2:���a1����%�d�*��_�C�0�87��+=-�=\�V �ԝ�#���3 �;��
J!�'�����o�J2[�ё8Ia���g��P�;P�	!|��������v@B�$��i���`�{�C�#�.:2��b���7�R�4��s�:��?�>��w�@�Av�� Q��/O�D#sS��<����_�$ LnN�CDL�%%�J%Ww L�(�M�%�H����S�Z�kq�?r� މ5ݚ=���A�%r�ъ���}�0��n`$���,���'�0����IƁ�u}�[ڹ4��9�)i76�ȸNPդ>he[ *[����N�?����w�ݦ} �5�L;p��,X�1F��ZtN��u�c1�pHX�������(/{�P�Y�2���^5B	���a�O0&u�G�_�3��I[���O�ۻ���$���"��ώ9��Xι��v˦�@3���r�kL�=��k|�ל��|�k �Oՙ��7_xDo�P�;��]��<({����3z<�N	�l@�%R'��ld� +Z~8m��MU˸ x]23���{��Kn�[.�be���o�.���8-�y>�|F��89��-L,F�GE"KQ����D�5��y��)�����.M|&7��:�ٗ�2]���2�+]Ǽh�B�y�<G��D����S���,��`�u�m�$�'��T/n�^�{"r���#y�B��WS�96U>zG}X9Q=�Z��"̇�%��;��=���w=���f�鈞�����0aƩ~:)��[�:f��
vkRK�E/�����nBB�vz���l�� d��@͚�d���x��ߞn���p�KB(���{��}>�)!T���U��O�Pj������d�����Ŭ�!ơ��O8R�GK���P�'e�F�%�a�^����z��e=�O�����д0��&�6���F\��A��>�2�p���C*!6P�H7�}�i�6�!;A���^xL�V�|��ͤI�������z�*����1o��rJ�}W*E%�g0��ˇ��F҃��k�^��;�X�X���i�Ik�,~s�DҺ5G�\0
	�s��M\L���2�'A��s��$��d�I��s��8��r���Zƚh��F_�`[��������b�K�����������E�UH�(C:��R��g�e�=�	�bҞ���H�嵬5־G�Hw�'�c��_9�FG�#��q
�1�z������7�&�ph^��#i8�&HۺyL�����p�3穅�+x	�zY��eJ�LW�Y�zDX9�B��\�Y S5t�6_��U1��E+"�)�P�ZJϥ��8`���7N��)�jwF�1�>G[,�������cT��D&�s��D�*.w�!�7��G��)�@�B�x���9}��e��'���B�f�6d���ݮ��_��c")_Ǣ'�`��[��!S�Db���^��C 7��rf�=��خ�{�j��PCӧ�C_�OU�� 9CQ�	��C���&6?���Ўi2쪰n`%�`eH�uo�۳%IY�����/��5:������=�0���Ł��7O%�ޢ1�2Zt�\.Cͤ�,�5�O��V��r�,��8t���C��y6��
f���Ń���/�H��=�|����r�a	Yѽ���ū�y������h��6�gU���4H��[�p�ƶ�[}q�Q�h�= �1�����=��!�6�SB�\�Ռ���{.t v��W/�^��
9��?k��%�r_�I�;K�Ը0�rh4�����v3��r�&�YG��h�C!�b���+Q\�����Ft���f�ِ�k�F�gT0��rFKG�ǏG�����\���wDZ��6"�R"�C��ي�L8^J�ץ.^.CrF��f���Z�z"�����o��Q1���3�8%?�  `���̶%m�*�+_(�]f� V�����5l�qy_E��0 �!���	A��v�dCz^ڮO��z��A	}�5��#������]s�������=�$E�ǎ��L49�tR���Ȧc!ϟE(O5�	Ƶ}�%E�����塗Q;X�A��]q�[|����;*������i��M,�~���8Yӎ��B����x_VK5s�4L���\@@]��E�%��]b��A{�M�׀r���}�5`�����ԑkS}�Y)�K!��ۯ������#y~!�*Ն�*v:�Ս� �fpg�Ѭۇ0�U�r�����l����y�gі9��wlT��xD�#�ʥ$� �M(��6�y�Ų�q�#�"���e��G:�H�ןJ��Uj���t���R�Wg���8o����ak���<�$ИZ0)aj�G����;X_%B0<�(t�0�-i�I&x�Dq���K��ॄ$�,�a��������[M� ~��!���\Vz�Rѧ! �����	��ɞ�L����|vV�&��(Cֿ���r(��u1p�s����w�~�gxB��d5t��-��d{�vuq[�jYW~��lKE�sה7�]���T̝sf�C�5�ȴ�n6p�7-�rQVW�*�2�$�+<��r���g��B�)��M��#(Lܪ�/K������G=��>t~�����W� Ou~g�L�)��3�U�ݷϰ醰
��r'dIC�HzΔ:z��.:�C^؝����h�M��G�mG�3]m�y
�u����}A;��e��#��)!�M�tRr	�1T]Z;�������>`�2�{c�D�l��m�%ыwSi��e�DN��;�t�I07r����i��{��)�`p��ETqua����v�67;5#��UC0�~l�Y�@pdRvl�͕���dT��O��j�	�L�b�]";+&uS��܌���',�*��Z�ӳ+�E@�X4�B�٢(�H��ׇ`�J�4��z�I�x$�_rh�M$lH�T8�Ԥ^�ek,L���%��5��/�(&���]l�#=ԟ�x�t|��2�9||�@����,2{�ז� TO��F���[�e�5�Τ2M�l�}#���c�gּ{<z�#�'١�Bޫ����_&���.0�'���P�4!�P�'*v$�(�Gsޔ#v��p3��Ոs7_��F?���e��-�R�O{�Ya�_�����{HcLK_`#�?Ҁu@���mx+�s��~��yϚ~/��h��7������G	?�4Y>m�*�=?�_"S�T��"�}����,'C��vW�V���]�������]X���	�\x4��hlN�D������E�Ѥ���қ��ljR�6J��n���*�d�❕��!�1�|!��_-�;�jMע�TS8&�!x���*a�������|���+ܸ��{"�g�8!�E~���ܠ\��2��K���	��;b#�����t�02>�^#�.�t�1��&�tZTڋb���M��*�J���Kٵ��,|�wT�!�8ٻq�	0��s��`���a�~��/|��آ{�������a���m^t���)��8h̘�_N�M�-�v2g�3��<l�������߈�0��"Or���9�
�xL���^*1����*z��q��mθUҲ/7]��,f�{?���p)�J#�c� ̘�n/�T_B;D4���mC&ș��� X>7o���Y|:`\9J��B�^%E̵���.�0's<2ҷ ���pn�\��%�X���ʡ��I��A�vHi\%=�ݳ�,ڼ {˝������|�WE3`)/Ur�-?MC�d�[�E2�
����@�b��4"��+%�Hu-�{���˵ԙ&@4ͽ�-������x!/�H�4	��4E����B�����QS��a_��P9��N��E��+�����[w�֒�1	�Mأ�� �xm�N�)c� @jy������ӵ�����\g�B�Ȳ\��n:�d%�+_n��	Vh9KQr�e�ƺaEQ��1��er�Yk샘�~K�?����'��q}�/��L�oa����S��@/��*'o��21]���/Ä#�<��V�'��f�%ag^�"����n5�/�?&6Q1�T{�.�0�B7t3�/2>��N�|z��ッ�4�)\K�������k�׌�k��m�/�k�{�i��9�̃=�,.�~a���b�j��p,;;wYdy�����f�l��yn�X�>|�;=�����.��Ι!t�hD	,���JǼ�a�8��vCuP��[e/���ި�������S��-O-҇�\Iz2n�O�čDqG� �!i�dؾB�([�������ٺ����Q�hY�nd�f���!Q�lI����
$M�%�O ��>w�In�t��*	��a�������n@���;��dG��4�)+-�<�C��F�}�v�X�\�x��bڨ�4$�2!�����'�!C�_x?O�6Ag�G~ӳ� ZF����a?�to
W~)gsh� ��$܎na,@��u�1��n e���=��z{��4�SQē,��'3�Ї���e�|ɦ��'o(�؜�6����K��Ρ�����k� #�4�Qb��E_��Q����\	�5��� (�;�?�+-w�X���9Z��&	�͠L�p��!�����4�E�R�f�B��|��J�ۓ�°��%��V�{�n�W�a�M ;�h^�z���*�"s?��h�Z�/��W}n���!�VD;K)$�U�1ؠ����p:ZT�I����uJ𨡐EiU~zaC���ɾ�^�b��(3�4����l�#'$���{J2�8��IAca���:��v"�Et�xP�.t�P���d�8�Eht��ɩ��3;�_�k^�9�����l����O8)+���1����c��������Ɓ�e_5ʔ�EN�P}�D�����@�߇i鏢ߎp�0|�AX����v0F�@{JI�Y���!LX/��&��$a�N���qo2<�`����]ŕ#{'�ǂ}��>[�J�Q_�XM5�e6���)����� 1H?`���Hk�e�u�pl�Wu�v��SF�n���H�.�0.�9��~}�0A�ۇ��B�{��i�EE�)Üw�V�e'uJ�����~>�D�,E���0�7=U������ΙZ��P��}*�9��������p��[��i��˒�,C���n]5��*eK���F���8 $\�Q��{�BZ��)[�c���vˠ܃��-q�h/�4|�I:�kU�`�5k˳��33#�;�$��m_�dW:E�����[aS��i���s�}_x��������?g�
zl�H�B�^SNSd��
Wh��gU�%�G�x�"�+J<�V:����s�l�?B�|�I �5�Y)�L�$}6����!e񗅝�cێ���q$8���Άrdr;����3Sd��  �Lb�R� �����
�[,�nUWA�7���+.���˺��Hs;'D�<S�wJ��}"9�7��Yr�AYʳ!��i���u�Y����a ��T�eG@OҬOQĆEX��.o�v�6��pρ!�+y�G��=�������7>�B�z˞=T,-�w~m|҄]����<�9�H�*3l���0q���P���x&���q�:��h��ʥ��k�J�N������+����}4��������Za�`���3md5�3�d�4��c��St�����&�7?��qa����CP�S�/�U�����ؙh�Tn��P��7i�k��'?����~iY�m0x��gO_��5[K�:�e. y\��΍!�q��~Й:� �v�"]�"���/�G������e8�IP��Ý��j����;�2tIE���=R�V�@�@3����`! �/�N%Ki7p<\���2$(�Q��ʤ�H?��k���;�o�_�߹:�mDyף��Pp��[�o	r�p�9��}����>�G7P*,0��P��Gv�@�����|�} ��s��
�NnBgZ��� ��k�CUO��T�d �\��$�Xx����\|�*�r�wb,y��]�G�~�HQ�a:щ�x\�@�Ɉ�l�0r��v�&	�xT?�c�	��<��T&�U�h��ٵ�%��T=8�-=�5���*
eˮY�"�%��$|q��.�/��C�g�oR�r${�!9.-#vn���F
.~�%$|�[��,ط��2�� 0O��I*A/R[�P���(��\�h���YV��C��m�26Өjۅ7U��<tɵ�:�șx�AOplF��Z�wp@�u$��K`��I'��6�Բj,lR��]7!>"�M�,�B�O��tˇ(��F�K�>Ɵ�};�±���#F.�k*� ā�-a�<�#�Uh�E��m�CExHEг�S���(j��:�k�#bl�@'�E.��)����a�fnCyzh��)�;����m��T�W�V�m�rI41���X7�;�/�N�	[�<s����C�`�Y9Cא���X������/�_��%Ձ�������O��#(��SH���'&/]���M4�����E�i,�!uNT��7��;��-��"�gi��i��ouz���f��{q�խ����>[K/�>3��?�O�k��<�͓󾏤�CD�Ͽ�wr"�u��Mm����	V˅��r	�w�p����N�ҳ��y8�&����8���Y�8PB&��E��VB�Rf-� ��7���l�J,�u=��uvC����,T�t���S5���%���N�'C�}��]��oؠ��_�֥����t-����<{@]<C��H20���:�[��x�wA��w00����,cF�+5�dB�u��ڜ=��r9��?�%�;0�Y�{8h,����f�듸��l���ῳ��h��o3<�ȅ���Q@zNX����U�~@z�	'}�1N4�I���(Hy����� J���Bk(Ҵ�.��_�E����p9p�%?�p�\r�~)�\	�AAf�MOQL=�r:������}G�LB)�~N]����k[���O��W��RL	*��<J���1D�.)�Q��}�M!�5��C?��QK6'u�� �����
, �ŊI��^g�z���;F�e�0�� t�Wd�h(��;�.��y���택�u� EN��Yߢ	K*�^�VB6�5���W.�2���.;-B����{��[�u >�rzʓ�V��$"+�0\]�вX�A�Xiq|R��عy�oѣ��l�M�N�Ѕެ2��F�e�t��a�}���En���Ν��ĝ8@��j6}���<�����D�]��1��
�d&E�K�)$�p�M���>+�
�V�=�d�y�$�ke56uPq�S{:���9�)[��Y(�t�	�������jM�E|��(;Y2ռj8h��,�!i���z����cr(�j����d��R�)���t~�� /7�Đp�+���}g^�7��f��A�}��%E�B~�<ᥳOT��hb#�|:!�����ɏ��	fmG�G�z%�:<��J;Mϖ|�*���.�R?V�|XL�uߚjє�~��]}��rY����ڀ��<,���Q���Ú֗T$@��'�B��[|�R�`&��
5�J���a���"�{�_�HtD2*DY6�os(x������5<��]�g�!Ğ�Ga��$_��Uju(.���'t<]9�\Z (���z����oܘ�վj/�.r��8Pu�3������\��ޕ�x�R�ٞ\1�o(��
�#%��{�5}o�J�c�"SU���2��%N	��tO�i;�	��\Dό@-�H��*wbK�P��S�Y\%�d��ߎ����2���|O�+F��������7��R����ǔpK��v\�mC3�2�C� ��rk�B��:�X�=�~�u�}>U���ZV�y��"P���_���z�F���ս�'���S��na7;F�6i�_���ͤUFE��V%�O{�u�Rm��9#z{�o�\6�����L�O��exjmD�����
����/b�:I�*��������lԽ���-tV�k"T���\�4�.�'��z�e�a����ޗ � 1�f��55ր�����=;�����Q��'�Շ���{�Hj,n!���B 2q}���^����)����E
_c���S���w�qʙ�w��)�IG�Al�yl��2 ��T͵�"o����ev͎��l�����1�cb�lH�\q4_��������������{z$>�QC�%����@+�eh�'^W-��?��<]��#Jd<�]�1�*�#�lG0��������pqa�g�]���#I�U�Q��P�����ʐ��;�vhb�sh�Bȳ/��4Xrgm�[A|��\��2� �H����#c��^Yg?�U�V���h��	���k�H�
�_.��8�D�TQāl���[�^����� 1����a����#���Ñl�n#6^����:Zۍ���Q���NF����&p�5�A�81���町�qRP��x���+�ÿj���i�7 2U�0�sy�=���F��� ��p` G_	��$��w�����l��I����pLZ��,S�n8Ge[k#���ѷ�c'��^4����3��;
�V-w�wʱE��V�w���݉/c�p��	��p.ӽ���(�9gк"
�������z���<R���{� ܃�����y�R���
G���F���z��4E�Z?�B�8Ni<��� ׯ���_�0����&�d��RD��ɮ5d'��x�H^5�����x@M��/Y����C� ��V'�l���2T���"�~G�g@���dh������TWF�d�["n-�b���olvn�X�9U��x�SRu��}�X�V7v6��ܚ���I��$�*Z�L8��t�{�  ��N�4	���M���.-��0ׅ.c�~����)�8CĒ��Uľ��.���~��R_#��m�'��g�$�bC���ϱy��>ܤ��`����m���z��`d���p.��=�g~�4$����0�#�����Z��p��M�0�\n7>����ѯ|�bð4I$�߻\�xuH`H���H��W�`�>xJ��a�6hR̝@���NY+9F�x�%�D��@�=F�c37M#ͫ̕"~�.i���ַ���A��mС��Y���դ���a"��
uN�I�f�i�fN� x���O�w���Q�m���wM�cQ[�(��Ȭ��UZJ�h����Bc�e*/R}�-U+������)'a���l�G����ɕ�u5P(�d�?�y1�.���(w�ʾ%�V�&��A�⮙�fm��݆���gP�6֞*c�pk��Ek���������6P���a�����T���� ze���k��5��RB��L@ �����
(�vjuHźPn��!�#vޞ��	�W�k���,���/X����8��@�$�?*�Z 97��ճ�	���ۻ%\C�fz�� 1ٲ�5E��GcVP�/���Lk܎�8a��Z�fy�έ�\W/u>���#.p݅��jr��d�)�tm	��("7A�&R�����RX��'	V+�R-�2F�|��,����n�O����#e��3�;3Nw�=�_�$�8����y�~��e�K�N���R�Y�=����!����P����NY9~������O�j&	�<h,���e�02�lV�w"- "HM$~�+�/����$��B���6��V��@��!����K��n;�E��!::���U����ےI(7� '
�h�;+B�$�L�����
���@���5��{�����~�:dG���xR�o"�#���}��3,�����'������<9�Hǡ*y�{�H�]����_��Y��u/�@Ǟ!�ݼ6��֪�������V00)g����	nT,�~藱�ROj��g���$Ol]�����D�����}1% RF�I��
���e㘟nF��6C��}pV��xl���!]�������v�[��s ~7+���4�W58�u���X�m�NW�k�V�}ܴx����A5[qdy�H�ݑj��о��R}��Z�~������)8��7�r8^�L2���X��ཡ�g]).�`k�$|�r��a&����:ο�H��t�R�;���6 W��/�ͬ��Kn$]�H�G�#���Z(�u�Nگ��p�`��N)o�53�f��X8Я�r%���%&�<�'�S���Pc]v��X�3!�����^y�יw�N(K��ˈlO����J�kO�7�R��mT���{�� �f��]�����d�<��(]�8�i6CzW�ő/ϲ�01s/=T��g�~�,.%���"{�h�5�Ji Լ}U���{��aj�c ���<�{�8"�3Ɛ�8�������.����1�Ñ�x,'t~x��BA8����3��:���������vbp��I%d']�I�S�!l�񏙱#�/楧2���L��~ �\D��ŧ�L��հR���DR*
�<��˳�b�<q扙���֒Hh��H"��,�_�m�I(He\���=�ޢ�.g�
�{�Q�3�v`��6�J��):ߏ��y�� z�ZkX0B�[{06'��E?=� ֿ�Z�/	Lۺ�
��YH֏t5,n�I	��_��r��I��ZvٗR�E��e���?��n�q��\�֝m���E�\r�VЉF*ߙWṵU���-?��C��	T�I\��r��g�FU�gF��H?��XC�y��ә���X�AS�礲����}�]D��EK�?��r��$?�5)VH����^LH�5�2��&Z�uR�C_5�P~١yU��@�3�o��65eN8�8ʕ����k���ޤ���; N�;YRВO��O�ĈCC3�S�]��D���rݚ�w�庖ƈ�\�����'�������f� A*k�*��A[��5�x�����Z����y�paQVE�ߝve[/��!
�3����p}�גC�k�ZΝl[1 �rؕˡo�BG�a�}����11��s�5����9����дx��Y��(� �=L�;�*��˲����U�p#��g�����K�V^;	
�H�ձm� Ìء*?���z��zL[�D���0�1�`Q��w��{҂�*
�ҫr�$jӉAL���^������4;�q�}2��6���Z�L���eW�T��T�O}^pv���up�Zn?�'��^���JǱ	`w��s�qV�Qq�	���������fd�6rf�z��ѥ��I=����t���\\.F��FW�>��0��ϔL��XT�i(�IY�ѭ!����%m���ga����cY3�p�k�X��̡����p�d�����%l��T5��pyDSD;����J憌���y�:]L/�%����Wj��ż��!��PRj�"4o��mS:n1k^&׵���+�����D��鰪k��hd�4<�B��6�X��P�1&�*�fX�����lk�*e/��T�~sǽ�U���ܷ����AS&���"�J��Hap�6|dc�>�Z���!y��
��,��x}��v��em���0�H2��a K�7��<zY���b�$��6ᔨ��<G���s֜�D+���+}�zC�����J{ �ǝ�0F9_ǟR5�Iy�ey� _?`��O� ޖ�#������p_�,N=�:���g|�gAG����=s�G��7^PEs��G��[��_���+�'��UJ�;΁��?Q�La�ןV�"��p�T���c����RȜ����9	�Ul8��6�.0�
�̡S�
Cr��6<�r2�����ѻ�+h�՟�e�|�-�6n�ֽٛ˗D����Vg�V�}��Hnf��_���[	"TI?���܎`[9ܳ�)ֶ۬#8@�Q?�ǵA�����ZgS�N9�@t��.�O9V$��*6L)vw4��--phS����ȃ�-:��@�"q�:r�n��xe�(��.�C�����������sj�%Z���m����M��[��ĭ��v��*wj�G�^YD��#)nx�v�!!�3|�(�ۤ4[e1&]*��Nt�6�����Z�d(�ǁq4w���������@1+MQ/ߛ���T�?/�ơ|An�WZy]��^�5�Ϥ�Q�e�[j��q����,�0��,��m��)�*��
N���<�Ld�gp�:��ĺq�� �����{��)�-�@��һ�+��*�1����$1� h(��~6��!�+^�]Z��XAK�ʉ�^����ɗ'W.V����*��4/ Wg��w���L�<a �f�J�y`7u��ل�'��2y.R��2�3�~�����ކA�����}�s�c~��as��9���Z����|(qk��ry�C��H?Xn���UI��8��ݨ2��,�%0%�����2�OѦc���d���Q��~�z�f8@�j��e�� ��&�г�Z�jd �װh�j�4�w�T�	P�S��m�:2�]P�$��1��f��c��Q� ��P;���b�4K7<�i�8���eKL� v~�l/��76�h���#0R��'Ŧ�H`�[��H(�t|�V�GZ��EQ���20�M>V���%���8['��h=/��Ć���E��/L�v��3cǽǡ����/��@��o�D	�w_=K�K
D/x�;%2�&�l��M��
����a��5��[8i�?��;�P�����8�	e���(27��7��ύ��t�.j�β�(�ƅ�LIe�x��:V�]B,Şs�P�Þ%�k$*�sX�P�L���7HJ0�w�䶁� Uz�{��b�!E+֒�nc���Uwm[Y71��~��4.xE?���e(�+ֱ�dϓ5W�4��@,�*or�(|���zV-��w�[�ը�Ń�����Y{�-Uvs�+4����� �W����a��Y��p�RF'�Sq�h�r:S��)��s��u�s�o�/6,RwlJMt2� H�w?@'�K�#�����f�i���\�!.i�t�����t4�C^�A�
����)�")���^!�̡4ޱ(�G8�9c�7���
@kX��0��E�	aˡ	�� ���:h�u��z�A��a��Jh�D����V_F#��#l�O�=�U����і�e \K����_7��3��
�1H#CI��WSU��Fξ̷��{y�D�*w�!e�~k���o��ÞHZo�xƊ���/z�O.��?B�i��djgpn��x5\^�.U[f]��s�������+�4(����<B�j�GP�X	�*FQ�x}7*d��ʛI�*���D�1�Z�w�	ܽ����pZd}@�eN�k���2�<�{����*;:6�� Ԣs�o�s)�R��0i8�e|��A	 ��)0\-"t���U�S��.t]���oǗ���������c��"'Kl?�`4{�q_Ǚq�x�#���6BV4h��~��ϯL�Y��m��cɕ�m&5�N�
�/�ꠅu�L�3���8UBF_#Pz7��L�Kq��Ӂ��,w����;:�`k�B���3d��P������!�|AV.<�����*#�H��H��{
�Uh��.ynz�Q�����}͡��}ZcT�Y&�@Ԟ4�%���iE*��,���%y���Hk��JSm�����=5$OL�gyM�����π�s��ڿ��Q	[�'g�]>C�2�&��:9�Eϐ������-�ۡ�:f�Q��3tdB>J2� ���i7u��Iq�]2
� �i�;>��A)��p����'-&�"b`iǉj'�'؟�#*��pK!lb�����W�<�@���ơ]P^H��q3�m&B��|!	���@|��F��3�͇S$o������O�� %�� #@#��n$.(	:r�c������U�!�"�FI��G6��!	��@���3��OҶ�,��쁱��,L���0]zO���l��&P����D>8�TF�2{S[�~g�y|���Q+�hИ]`*e:�wYM��hfv$�J�P)*t)r�Vu�񄉦�Y�,-��^�C�Mn<�b�zS�:j������p �[i��E��r,���(�"s3N��9��������{ ��q���N׊��̵HΘpp����3D'�������o���K/�S�.87`��Kx���K�6s���Oޣ�!�ڱ���U�m6��y��[��7��W�4&�Cqjeo�wϰ������v������0��D;�#/5Sw
���H��oAp]¦�qg$�?*��G�Z��� Si9�m{���O�yO�<L��;Y��e�y��ug)��'VK�Qh�{f��5��m��fk9�mXk��^1'[�x^d���n8�]��o�����9B,d6��~o+;/�KW�1���y���
�w��9E#ؾaf��l�韻����$w`�޷#�J�����t`oe@1Y1�/�C7 ;�w��r�,K����6I�~��|�*7-����\k=��װ}ؐ�$I�j�'�˜�[9T�3��
A=k��n�r���T�~N�e8����4�_���=��yy^�!E�L���P\W���U�"J��MD�Hïzr�yQ��CDah���y]K���>���n�F�s�bh6P�I�!ZAS�g����x�
����Y�K���K��#�fT4V0�k���?���fVc�x�	Vӳ���xkX>Ն��v@����ǐh�%��г��3�����f�A�R���@�`&�)j�����)�$x�S���w�\�?)&�_��@71� gym�ԋp��Tc�7�_����ۄ1�s6�V�XB 36�af�(��5��eAD�J�"����:q5��x^�(��;��@�����Υ�Z��VP ��2M���.	w�e���[���2���O`5f�aB������F_
l�*y��k���6�`p�� %���<>]�n#!M���DI�<C�S7�{]��E+nn��f�@r������`���d�s�$�?Mݝ�h3�5�<Y|�E���Kv5}'�C? 3�}�S��^i�"RG���R];�[F���?F"-\,�ꎍ�� '��B���K��6�vb�ڳ�B�bVH��ˁ�=��j`ᜮ�ѭ�:Ӥ�N��'ڎ�zО�>	�C6�z0��G�����`������*��K}��G��E�n��2�\n���ٱf��e�M6۠�1�J�4�I���]���42��y���5SF%�m:�ˢ���K�R��<���~�]��|:Tg�(�������g{�!��o1|��X�M�_)�`6߫0_�d�<*~)����Uo��K%��\;�S2Ĝ��5�'uR H
@=.�YK6Mz=��A���h�!��Y����J�~t�����$��.y�l�[��% �\\�=Jb�m��k""Vvؙ ��C�3��9	����F����E��.|U�[p���ګ�)�<�i#�!���B�����H����X����V���3����_���c�]�^������	�eU\�Qf�a}� �u�E���Y�u���a�9��f����<�5b�	��V�^z�V^����LVm���s�P �jUO�ο������g�N�%�u�*꓃�4e�h!,[ �>=���zl�����>/���Gh�"��-T���ʮ���>���}R�E��W�����2�X�hD{�Lr�=��U�*���$I|By��TP^�)����('�X��j�_F��?>fm@ F��V��wOwy���0��=�T�Q�)��� �xi�]a)[�ίW�`t��`#�^�c��A��R�!x:Q�Z��Ej])1���Gk�=��Y �_f����|sQ�gb��*>
Տr�D7A�t��x�l����2Y���Q��ڗ�,���<���l��]�Go���{�ݐ�]r�c�
�N�q���!~[W� �*�a��Բ/t��R�1�x h�R=�Ӧٗ���:H�
��ܝ��@���2��F*��s��*�q1Tr���C̉�.G�f�{J���vi� M�9Qՙ=Ϸ��iDћ���R�g{5y`΅����L���r6c���@?��fm�
b�������b�>> "<�Y24R!źV`z�81o
�f��X)�K�ʵx����i���p��F(����h§����;�,F�/��Ӛu���,�@��3�q�����E���$�e4��Q�8M�,Ia�_�sU �� s�/z+#3�f�y̸�*�ҋo#�W���'n�О�d��3ӳ{���t'�9�����K>�����]�F�%�`�#>4��!�{�? ����Cԩ{Wx��k�:��$���t�\:���~:'*Δ�މ�D
�\�	�43`����Uj��ϫ�9�	�+Q�?�-6O�TW-�~�,X�g��.���[�ɭ�
�T���^r������F��n �ƌ���dh�U	��q���@������/�6�D�Lf�y N�;.YTd�Y���>�2�`���`���$�V��E�.���T�Pl*��[�xCHZ�^Z{#�b�����/D�0I�!$R���N�d��輒Π\�*}A�$�_c2UM��s< ��\IV��ȢRv�۞���D�j@亙���K�X\d���N��O�˓�yU��TM"�o�3������m��*M���Kr�kf�Ҝ�|]����(�,�Q��ƞQX��6�''�;hڋ���/|��̋�r������+�cJ��6Q�[�<[i�~�'��m�W��~0��r^��n$���8��=rC1��P��BR�[��b`�&��ڞK����RM>7����41$e��4+�� ��R|��q��rJIAX8��S�nc�D/?���ԟt���t�{V�'��,�� �ׅWMP��IX���݊���ם��(7s�����U�r���v��E�-%��7�(�Sj��k�n���~�30�>������"��V��إ"�����B?���x��`��d&nE���lvi�_��|�@JW`RU[�q��0�,e�烀��Y�k �(�*�,��Z'G�SզI���;��)]rF��5�Wȣa��Z�nVt6�_)�����ޟٚ�>�av
;��2ݞ>~=��STު!��oq��)/9�X`���q�7>�x�ro� �Ҡ�_D�cz�$�7�)_=�����,��1y���~��/g��
����[ �|-1p��,TN��K�\cu�����ΧIq�eC�$�.j3s6����f����,��<$ZT�s�=�
��?��}��*�
�o��~[��p�ԡW�� ì����oM�Z�uQ��;�����@����L�MA��	�re'� Ġ�.vS�my�5�����[<� dε��e�cy;����`�{#"�_<�(��=����85k���I���F�H�ӧЯ����o�q���F<����`
�����@��{I��͈ɀ����.m��N�!gOD�I��E��k�9i%�!�O)���|����8t��������3������^0�㮊Ee��)��׫T�	�
���e��t�?�#��������){������ح��*���b7xn�<����{���|�K�r����M�<5�rnu�ְ��1t��.����f���#	��R�
�I:�VŮm���y���jo� Wr�}�70e��Qj��w�j�8ёx_����þ/�ɻ���(JL�`�[4��)&d���B�W�Y�ig�z%��]8���vR�|�갈��y'�9ꏔ�Vz�<�w���%+K��ҿt�8��6�l$���jC/\&0�}��#rU ��f���_DNڃ����m�s|�J|7%4�����r�c�F�����R����$� ������R�w�b��eDh#���g�/�V
8��WjN����� ��d9��E�ѥ��w0}ۈ8���f�ʙ� ��š4�'ݯ�~������s)X
%�G��8�썅 ��?�*�\ͤqjՆM�{y���4S*�}>����Ox����8@��&)C��Qc��h!�T�hf�[� �ڶ���y�8��qC�UK����r���q�\�U��:iж��W/zu� {K�Y�҂P�	T�n�
���>���'��Zօ��ZgN>�4�.˴>u���oġ��oD�� �k��� ��:��'�{x	t��!�]Wq������[�fhÇ���w4c'�ZN���W��܌[�f@o�ʊ�*+��h]�i�.�<ا.b}	q�'�˔Giͮ< k��8�>XD���9�"���ʫPwa̖}Fo%��o�g��T�-e �f~|���y^�$"&��חY(�WT&!�X
$!������Yf ��������撒·h�?�=�;~ �f{̐�g�1b�_N�!q�O��o�CpV���s�D�l�A�Wi�K�O�|��+�(�+�6�g�]^?iB�$k���}]��'8H�I{�OF��O���	�Pm�I�C�7xob����]K���+�"4�xa��[�i� ��Ʈ�_��� �E�e��R� ���оL�
�Љ*+dIj�#�ŀ�ǀi�5;�
�˹�<�`>�o�-zK{y%� �������M��4��ӟ�j�>�@a�����O~$��k�8ӿ�٫�E�������[�S��.,�D B��$�&O�8΋5�Z��U�Ѽ�����m���}��FE,�O)E�$�v������m	Qa���Uu�ٷ#��X�g9�
��kf})ZQo@���ڏ}O>��H؁`Jy���S+[E�ҬxbKv7���纬�w��{���_j4��!��p7GO$�t(��X<Mj{�o�L��/Z2��b�T���l���F*��)sӤ0~s�d��?/&R��:x��4C- AJ���Ze����U���񀋗<���Hmz׷?lF_2�_'t)���N�
1��g�H��e�T`9c��H�VG'8re`�8����#��P��������G_Ε�[�_*	T*'�˷U�����c�(l���S��*;7� k�@�|��d�# k�������U���\�]���uY�ɾ�ZUg��B7�ė ����|`��=�t�l#���)EP��v���pͼ����B	$��e�h����I�jc*��3��b�� ���R���.r�S&��0���S=8�� d'��k(�2�`0�/�-X%U�__�@��K���,LK�b�ήM.쬽o����'���r�]p�����VD�c��WA{eo{����Ő���w�-�e[������,'�&���ݢ��ʻ�ŁU������1/��˨�e�� }��M�ډ�ן����ᷗ�f�:�d+$��Ios]C�"T�W�>QT;��n�I�t8̄bZr9a:�:�p�����#pN%�:�!�a#�:8:�B�ă�JC������n��������y��ִI�'��-���	��կ�7-9���C��Q�&v1;1C<Ҧfb+B����w+�	�{mTe�d���̽��b��W{Yq���G�ȖZ�G�V��7]g��>�0�:׊�︾O��Uq��8q��Ĭ�v���+Lz�X<^3��쓤�Nkf�Տ��t�x�>4,ao�P ׎`�,;_7׏@ݕ��1Y2?��Y�Ax4��P]����7'Sh���[34b�̩g�j�����^X����'��A/�m���W���N��$�Wap��-����c�a�����\��J�;�z&'_������zc�"�y1*DQRb�Q��z�M��+M佡{�K튄���\ӂI�,__�oӇO<elR"�p�g��W��U1��P�`� �= 7LZ��|�f]�E�]X��b �PS��1�% ��N�/���Q��̰�Ƿ��8��4d�J���7�ZQ���(�.Xa���eռ�%q�����[)���f5�@+�~�XEɰ���j��-A�]�W�>���m`�Es�Rк�Q
Fon!b��8MX����ڣ���Kg.V���z����(z�lj�Y ww}knj��%�X�\t8k�Z��W^B �������/���¤����ć��� V��CQ�^M�0���H���H����T�?.�x�W�Ew�����bu:�;�~�f��飷�Uh��Y]zR(38+���H�pyw��QGS4��A�����$�Qo�.;�9�T;�!�_a+���ׄ]B�u�YT'���Bn���u;t�s3����D����ː�s#�=Ĩ0]��J�4�`����0���#[��o�*�U@dܫ=:���O����P5|T��t�^��ը!�������থ�f�+����sd�����V�!��d�9rR�Q�`�X���(Pk�f��q�c��R���:S3>G�>7�7��}!�8?>�Q�	�l�CjFo�ކc8�Ī�ŵ��J��gH�Y%:,�ai�����k���촄$ԯ��3����& ���<q���a}���⃑%����y*� /Ꮷi�-�#�	ƃ�{j$
�E�J�Ko���r%���D��gL�[�J/�F=����ݵ+��>�/x�ف8�=��+�? �cݬ��X�	�i.r#�D��x��!r��:�t`�ة�ȼ�A�)i�[�NU��&y�J*��RP��Y.�?�]����>��+�S�7��Cҋ ��TeKI�y��x��y6̵&_{1�ϭyIIN�W�,r+f�:�D�����s�SL$gf򫍩�R.B<D��8F�4��Un�\�$�i:K�|�O:�@��� :�r�ֳ4%��Ӣ���K�7^�]_��p�[���j�R�RDC��v����i+��K���~؛��M���#�(]��P���=i�(���K��}���c0'�n�p�)�d�#)���}<�L��83�<[�>��dn������ɔ�u�Qv<�J��[J��s]���߹,���Lƥ$�c�(ژ��d���7LiP�n�Ur�$��Π��=OcRz�hL�꟮��6P������Ǌ-�n[%��D�*�OSx�?	���2��EB��YXQ*�v�
�(�������\�]�c+�M��9|
��(T/�,�Q���`>�e�h �����fBȌ�+�'Jk�����K3�)���q����S��g�DH?����m&�L�
������5G�}�XVzCx�{�.�e����UE���-%��gq���H��M�ęá�M�Ug��ɘ���H�K-
�U�h�q@G�a�́k��ʤ�*����=���lp�J<6a��_�g��:�h빶�J��8��|��̏zw'y?�Rn����G���7�1.�%�'^0j!��y����I�C.�,)rF?�z4�Bxr����0Z�KT��]l���W��r;��� �'U�7��Ń3o�)�V�ks��	WWj�C2��]����3U�G���9ס�8�	O_�'tV�"�p
��<,�T�\�8�W��:�v�Wi��.\`n;e�Ò�k�">�)���Ag�"A.G�$�Q�#���B;k.b0ph���7���t@r�C��Mrq<�vO �p^s	�B�v覽�rn
���E��[�(H�$5TN�yJ�L�'̙�+Q�SdѸ�l��p��2�1�D�D2ρ#8���ӕ��f!���ξ�k-a\��H~��Yb����{>?]���l�U�#�yyh<�ܝ��cKw��k}7�>���L��
]�����
�l�Ue�+�؊����$����MS����+����46�_�f���V)�nm;�- "(R�����^�D�h*p'>�O`tV*�1�;����O�y*�v�5{�+���i�.�0�DX�5�"{f���:��{����� *���H�y�Y��v��p��;��U�w#�N>�jwT�����8�sp����bI �c�4ZQ�s��V`�����P�܀EVSP;�X7�p4z�4,��l]A��vF/��bJ����;M�Vn����Bc��d����Ϩ�p6:}�te�cƟ�T��KG�����P���1y,��7�Ț.�����y}����Ҥ#{���T�&�Z�W%ԚW�͆��	�@�ru����h�pE��霍����}S��"���"�y����9�B�U�W��'p��X�H ӄ�|�^xt5��=�a��6���N���8 7ʋ���lf�펋Ͽ[`��i)�KPX�n͸)�)���b�P�?���ބ��%�|��|�	~�9��x�_yN���y���$}��2�g��]��֛Q)#>�:G${_y6d��t���v��C]aF�#������Y K����0��]�2��o2<Y���(U܊E�}Ue_)d裵0�`n����� qJ�v�L���o/��^[�4�*k�[��	�xm>i�Y>�Nw��m���kv���E�u�9�����C�8�(�j��IWW��&��ot�L�T�e�~�fV±;�m����2�ݨ�zg�L��5]\ X��4D�$�� ��\�B-��	��悌e��S�ZkCJ���8K
P;[ãw�4m���@�1�|�^{�Qp�����t��<Gmh�Y؁^� �eD�oev���zQ���dO�$9��e��c,�'YR\e�t��a��9;��4�F�f�w����ˮ�׵����]��s�w�
-��)���ণ~�J�H:��[�2�P��!>4:���ZKu��	z��5;��l7ZB�9�o�z��N����7{��Yo3p�p݉�^ ��i�F������^=?Jfw�-6S
/��G��B*�ґ���y��+=b��T�Uu�,I�b1�*G��x��n#���yWq6�^B1=��e�X=ˬmU��?���՚o�����ջk��r2(�o�, ��6�j~�D��.ִ����j���]�Qv#�d�s�^o(�v;�����S6!��:4Q�D�|�e^���Ԏ�Q
Rc���F�.Ro\�����u�%5�C�p-cV4m�;;n��Bx�o8gu"��+L0��S%)�0y��&�7��F#}a&O�}��=:����~�f_�G��ǫ�OF@������9��<�뙵�v����	O���j��$�k�V�V?O!���z�t��&�D��W3�6��:�N�c�����z�7�.�/��ա�Ñ�#��nOI�UƳ ��N:�ł���Y�ĳ8���b��Yj-a���!l�Zy(��J�.��S��Y؊��[��Vz)M��y�et5�l�9�.��=	��2�vd��d�����]�*�E�ٿ]�"�}�Յ�)��J����_�b1�/a�;���� tQ@n�#��1(��H������N=�M�J�����PU���vCs��ϊI�p��Z-���n@(�o�Qj�ʵ�S�%G���u<p��������</���swi�q? O"���&�GdR}*��� ��i�M��<��&�=4��@d/[ckbI-B>�O�YD�k���dN�4�A����%����"4����ͦ�88��^~z4l�y��'�������s���G�#E,y�.nN
L4�6hI� �^k�#����՞ ?&�M�0�U*;�,��NB��l�AŜ�B��&C�(k�h�ؘ?s��,v���CG�jm���vW���[��Z�_/c�,�K1>����-�t������g��h����$t�D�l�\��`�5 5�Y�f��|���	^��*@�%�SD�$���:d���!��7V�$�}�~�3j�'���.@���R�G�)��R���E�C��뀈�fS�_SZe�4�5��lQ+�
k�qd��E���o�ko��Nk��dTD��ِ�y���jKo����C�}!%����Y�0�����Bz;s�z=W��=������sVc���3�e&Y�$W4�A�h����5���Oo=�n�ut���٨��ߜ�q[�~���ݽ�_x)�EH����'[6�N�M��m�{@{���ߍO(#
�����ӬUL�J �v�qKCtr�������K�z7}C�)>Wv��#B�tI���C�g���,�>��\��&ϥ����>�& �;�Rz��e���uJx�==��4ɍrX��,«0>�Q%IP���\���E�C�!
G�La�$N�Q��)�k���
߄�;����D��>J�����́�"m2t�WQ"��9Pv���2��@�׿���`�cQ�Q�Z
~��%<�\����5ΡvC���#�6��>x�t�{2:��ɥ���Ш��7�sE���6��}���H֐�	:���Q��vu~���X6&"��K$c�Up;�Rو��ުiCT< $#���iy�:2�rzo���n����z�N��qh�!l�g5r:3�a�E�tV�+e����׼(j��;����ƮVL��$�'f��V����P��G� t-��5�]u]"�z�W�~E�!�5	�q!bFE�7 *��_��^�g�w_=�q9<�["W�SFa�����uC�~3k�a?�ӣ�Φ��fgA�\=쭐QtB��"jS�����~�`�F���k�;�����\�vܩ9XEq�.��Sa!Z�\��Gl�;܂]3�G��% ��M��ع!\���Ha,��&,P3 F(����2{�
w8��L�]�2.��;I�<��T.ЀT�v,�yx��p�Sd�Υ��p`�H���w$ױp P2�g�A���r����P�yՐ�Q}*΋��Y�VO1�)��
ƌ��:�Q��X���0�c�Y�=K�Q2�p�0�۴�`�(�Ҹ�@Q��n�����n�u�ܶ%�����]�H��,xm��7��'�����ۚM_����Ä{}��$o>,_���:�O���L�zC'=���Kd8�N�@b���k��6�7~�s�3���%��?�2k�Z*�����h|��kyc�_����]M�'B� _�1Վv�.,Pֳ�A��i&Q��_�#�����. 'RX�cv���o�Ki<��+78��
��o��t��:,�䨜L	'��&��%W�����v���]�w�4F��~#Y_W��۩"�`��}�D՗#ǂ(�&4r����o3ʒ���Z<q�����[_h��*��NĶ�~w���I��PrM�h�Ú��uu����LLw�tQ֣ig�0N��,�w4\����T�=U-�߹9��P����Hr#�Af�~j*�į~n�r%�v�@�����Q�S�q����x�;�#�<.�4�ea�u�XfR�uTF���r�K!��C��|n�d�ͪ��w!l@����o�^�5F�	���I=*�iѕ���������l���pOy��zV����D�ߤx{ḡl�w?.�Pp�	_-�H��:��k⇮�5hm���-e�J������{�X�e���-k>Αe�o蘜5���ON����#�s~!��_z"�+���W��ܟ��K�?�g����61�+����$�nj���"v	[�5
� �>U=���:Ou+�۵{qL����TWsW0I ������Y;���k!�����p8���1�G�TzPVB%0��VZ��!! �8m�/H�lxsfn��br'b\_i�cXW�c C�r��԰���q(Aʔ���`��./�,��>��I�Vl:���ߩ����tfj'���'�t���w�+5P�E�ꆡz�^Q#�z\�eE��:��ˠ���L��ų��NG��Q�$���L��qĥ2U���ç�$��V>��Ǫ�KIa�cA��#���k�i���o#P`��;?�>L�܁�+�OE�������g{:lrӥ��&�����4�����"�ٛ�SLB �G�p�_�lTk��Z�a?�V<}CVTbg�2�U���ޑ�2c�Nc�9���hB/�v:�����#��\�L�E诌�n�A�'����S�M'�q�	�����JS$a):e�l�Ej��b���߆�4A�gp��7���F�
p/�*��3�)��z��V|��Ź�6�8�"��ŚM�i3�.s�U�@0ԛ��|�
��$_ۥ��`�����~yf���5�Q&*G�t��Y[�J�XNW�X����N?ew�.AL���'H�#ɢ����А�Y�7��㠻m��י��Z�s%uN<]�����\ɬ�T�� &���n?GU5�/�u�%���K�){p�og]Fhb2%k�$4=�\@����7 ���C����}�3ql[A���V�p�g����ޘ������|PHh��=3d@[˛��ɞ�r�Y�l�����x�%u�������":��i��^jM�R#^�6T�_9���Y7ޖƎ�C�����t~�0��6�5������o�5vM��m�+�94���-q�O^�dr����ݻ��(��щ��k��3sz0��A��PsZ���U2�,j,�x��	tO]�Vn{I���ҏBܤ�p6����cH�D��J/�zSx<f��C�C>�?�yҪ���M:P~�ظǧ�(o�����sKקI���FH@�P���� ��7h�0�*vC���-����*3_��t�9�������lXL���J�2<���#KO�kҭ>O��||��7���X�`��۽'a#��8�oݱ���1u��7����!����,��2��&.9�T|��*�otU��ы��낺1K�^$&������+WG��l,I�d+���M��xM���O�KS��rr6S���`;3_G��C�g�/69���p�(R��-�< W��>ꈩh��@�%��Wk ��?\�
�LM�ã!��%x79[�M+�Gg^[�R����]�f����An+����y�򩝘�z|Xƕ}'t���g��M���6(�Q����=��4��Z��}�7H"�w�	�Fs��<�ܫLe]U!H�:���!�w�_�IFI�)��ս2���Ӆ��"�[��� C����E\�;'�����h�U�k)uQa�ؘ�~�7,e��S�R�w> �l�t��:����dڬ�X*���]�VЯ@��6U��>0��K���$!�X`�/��R�X�����!�aM�n��n�+,_�S�4.��4d��I�pAò�Jq����������}<���@Z��+����7�k���T�ԏT�u�
�j`������(`��Z�V�ђH\1�oUQG|�JPif����屮�kM\Nf@P	���0�$
����cxW Y��hC'�����p��+j�$�+�*�����;�L�Y���|��l���rɳib���=`%�=8(�R��ѳ���a:���J�=@ӆ�7�B���]�8R}��ZVip2�4�V�Ԥ�RXzw_�p	���u�}�g��Y�������wn>p:?ge���6`�D۟�&�'���I��Ʈ\�s>�T�=�%�w��S��V��(B��KDu��׿}3A/��+����UA���S<�{(X�|>1��Q�����J�=����ĕ�5JX�kr_w���n���	�=UoA�i�<�]+F=Lu�
��7%\��o s����Lv��������H��7��WE4��x�v�_�zx	zڈ٫v�5U�;mPW��/���2�_���ްZ�}�s��`�[�7��8M�w�x	�e�AM<(��ͤoޒEujg@��Z[X��0�Ť�Ѷ!���V�cIa�:aU�&Js�O2ܧ����
�f�~��K�9�?�Y]�D��Ľp�p��~7~�~�����{)�V���s$���,��ޫxQț9�6�^�Y��K+-~n׶�ԩM�|
;�k�$��#)�{��[G�C�czٝ�}�n�^��*�!c�3�Anj�N�\nҽJ������+��S%]D���JB�;I�xÑg����۳х���O�>�g>�h���@���$ia�W~��&AI�q��o���-���
\:��B���D��g�2�I�ɾ^j�x�e�ӎҔz�B͗����5��4��<�y��;���l�K+	��͍���d�n=���
�p�:��JѤ8��d�=�U4?vO��x��ډ@i'�1�G��Q���*��fJ�#=�b��^O�r;�I>�谼���"
�	��o?&�Gu�++�ϙ w�6F\8�DΌ�P���e���8��!�G�/�g�W��$���͢#�)$���Z������?^�S�J���<k�,:��b
ܱZ�rI�3�8�4]���D���~���H��ǖZ�R�U�Zk���{%�N��Ps25�9%�����wN�7�0��t��`z�c�"�kF4��h2�<k<����M�o���Y*m�iy�+��n�س���n3��SInRw(k�)7�1���u�����������nœ
��8!	�o�3�rB�/��j�'�8�f���Qm�����T�"L@f�[�אY��7���;Mb�~�}y�ř
W�L�/�΀�Eԃ�I[-�"hR��F�x}΅����^13���=�,&�q�����Z{JH�(�E�+�JF!���A��q����������tt�I^S���z���Bz}~�O ��H Ȗ�A��c�^X���p�������0���1bJ!�b1@R#u%�]�pA2&E��\	�zr2����>w)wͮ���.��~Q5/��|�}�j��8����O������-d=�V.5��6�e�(���\��jl�L5�����̄����|�>j���/��ɹX��\���?n�6�A�Λ]E��j��6,�[�5��ԥ"�}��+��vj�;E��
MCj��l��v���·�菼]p�����m�s){�������Z���@�C*ͱ�#�ɡ��e���-E�����%���]�٪?}����e�I �;�*ϥ��vn�=ނ) E�L�-�y�g�r~� o�2��{�/9B�'+';�1+��5��VP����;�����օ3ǃ:WH'�T������V(�|쐠$�Ix^`� �j�-��Wn�v��J�Z	�V�(,��
��hq����^6��v
U��'i, ���i��`<^�:��h#����sIk�-Lr,��2�� ��U�&:���� �A�zf�Q ����8]#�LQ~��oح|UB���L
��J�	��c�˾d�'u�q^� ���1�"�\L��U:�����-�_���D�:L�x��\	�`~H��BBS�7~ �DP�ٓH������!�Tj�OM�[]�]�Ƥuys�l&k_O2�+�řaf�)��>��lj���ȥ�L�l�(��EC��`�fM'��Z��6+arV.Q�~x�0�YDV��k��g�ڌ8n�3����P��D^�����|mswg*Jb��
ڙ�~�
��U��� ��1<`�J��m^�+�Xe���:�{��Zr��x~(P�p�-�td�#=�����U��x"Dքؐd�tbI|���ܿ��`������|�tP�\т0&����k�`�X,�2���{��� �k�L¾3ނ�<�}�9J�&�Nk-������S�#v�z���7G��V(��N��|�q~'l�vy㖦K��\P_-��ƿu1J� �%���K@@����6R�2@B���tS(d]�tG*���[c��p%dj��"Z*O�Y7�°�a�`����Q 'ʯ� ,^�e"�cDM"d�����30\��M���7�`���_[���|bp��5jU�kE���N�Y�)�R��d|��Fs�C[ �ʌ�'�(D�:s��%Y��|b�s"}��%�3�;�6H	���5���"= �YjB�`6�̨���W��
7�C)�H������:�Ү��Zhg�V���"�Ĝ������>mZ��m���ěǽZ��3�bZz��odg���X�����~���?���r�笫�ʘ51F��I�Ǔ���L�f"l��,�	G�p靵�X�`R��b�&|N_�O�i��%C�t|��Y�S]��_Wz�� NIA���^:!��ۡ+�L�v��τ��S�mE,}�G��"W3�<,�����y�Z�R�Pw�y�/w�;��N];0���}g��Y-��~�<���S*��ؽ#C�(Tp���d �����ϸ�S���B����l���k�q֗�smT�Sp�Xiԏ�T;��&��C;܅�$@\o��(#,9M�ˏ阔ƿ:�}��lsp`T�g��gv��
%ՉW�^̬��3T�?,*� �{��2H��觙 &��3 ��~�O{�D��
�s�2�SE������K�	D���4*ڙ��6s�F�é�%ve%g��8���pNف�#p�	�X�K��<�D5?�r>��eZ�6B+��-�$�I&ȻH�sPM���>�5�H�E,��0�?�ZC�|������a���3"1�%�| �x nq���1��;xD�����a��?�M��1�o�xs�ل�]�/�=dxo.����?T�h���4B#D������o"�[�V����w~yk:V;\�`&tty��
�m�BU�{y�$dm.g�������`�Y$pmls�! I�&�Q��QH�W��������K�-��Y�C���Ve.}dWY\�8�o�0���ڲ�ǥt��?]1�Nhi)��6�U���lD�I|OlõHI͋�%�G�˙��h� ��=(TZ�,=2��\�`DP��p��H�q3��y��P�f(_�yAڶ�\�:�mT��ě\�6K�G�L��{���1ڣG��",��{����3񈅓���x�|ۛ�:W��������6'��',D.�۫\���e�D���a�}%s}���<;�"�;��J�^�����7m����|g���'b��\����ƨ����N�6���T����B�p(RQX��X��ȶ{U��O����&�M)�jn�{���4���|1�� xob�ɍ���������@}�0E,��w7J�[�8l�+m�%����gk��ތA1�3r�OT(J|#C{8���.4�g�:L�	��5����2tӻ�Ma_�9ys��7 ��0�b��ݗe �-:��q�6����BdG)s�ߛ��vn��S�����ȣم��~C@&�G�f�ϓ���H��s|�n_����J5
�->ghZSJQ��n[W�p��ੵ�0�܁��ҕd���b	���T�������?�IC+k��_.
�NƱa#ѥҾ�΃j{ �.O͞G&�LK��%mi����y�����8�"���P*uA�dd� �̾&n\�*��&�K�������3�iW�����%M?�N���=�;�j�2�+$��:�4�xUJ��dY:R��`7۸IN���"3d@�4�ө�3��H}3��ΏD��rDz��*-D\Q,:���FrYt��E��h��6�<o���H�r��Lv��  �8�F��G<�+.C`�TG�mn-�픟�Y_뽇�/���adoq�Iԟn5+��5k!r�h�U��qN���`����/�h�3<���/�6���a���i�eyS���J.�� �{�=�Cf��f�/h�I'�SB6/8/	-(s5v<�����6�sյ���{�ϴV�@�Lұ�#��͉(u�msq�-s����_���U	�Y����#�7:�*a�V��J��]Q4�ji�y7��M;�$ ���Ζ>��[�#(����ݼ2�������0�m�xA���x�c'w:s*�Q�9pR�˸���V�͑�$�RB1V��u�U2ڪ`=�*٬čgㄽF���T��A���^"W�F~���xAy<��i�
�x�_�N��U�>3.�)gY�)��LFG�}���Eǟ��a�'
��#,MV��p.�1��W�\-�� ǔ�6�`�J|b�̛����@�(��������ʦ�AM#H���q/�^�=�7d]��N�'���ojz.2��<���1��2v�CL��<A�d�T�pɀ}?�<�}��+�>�Ϡ,^�œd���5����l�d?�n`�5��\LFK�[�1�(���5�����a
�+&I�!W⡬�XU�*_N��рs����D� V�Pxq?M�RuK���Z���5�t��l'�i?t�k��@��m	T��U:[����]��m���7_�댳���yf@Ȇ�<z�FYe���!����o��Y��*����4��'��&Ƒٿ�>]�(qz-������t3���g��>+\�����W߉�pM��v�$0�x��H)����!1�X�ui׃5��G��2au���<X����5�������ŋ��DJ' ��Ve2H�ȣ�n��� �(��p×j���U����D�&��u>�P`��u�fi���bEw,Z3�K��O����X�qE�Y�%���1�k A�|�fj K=��_4�SeFL+�u��Q�j
���+�J\75 N
-/Nd_��(�4��ߖ�v5t������}��ٖ��+yb�8-���'{�TΫ������\���.�%U7&f�`��جp�k���2+���5�����+��ӈ�|�G Eӟ����\�sB��F�N��DF�v�:�K._cз�J��Q]��._K���oű��Q7�y���
��G���Iu޷8M5�BkNW��u�� �d��MR�\Q��(��Ｚ�����ȕe��ߊ
=�<��/t������ �Ϧ5ִ�p`�]�}�̔��ctO�%k��a�((�27�@��ԧO�z�'�s���801���%����tP@k�� B}��:
�<Ңj}hL �I�%������Wm�V������gd���ʲ6��bu������GY����
�r�t���7ۯ�
$(7��H!S�������AR�-m�4wS���Z����T��$���,r�E�&bul�����gD��r�6Aˑ@�[�F�"۬�*V�C�ټj]�H��̩(>~�(»k����<��q���#�*	Y�����;���1���LT���E�6�id�{A���E�����S�aO�U؈|~dnB��G"=$����&y�7��q&�6��/̈�b[Lѡ�c�)�����r�����gl}�� ��K�[h�u� KU�)��3-�U����2i�Oy��Շ�����X��W���I�w��@T���:n�;�TD�+�\��<�������$e�^��ǿ����6���o�P~`��[�8
�d`����;h�Nm�t��Uk��=>��~4���gj��6�����o�%�ť�z^v�o�ª5ƖH�SM#�����Qm�D������Z�������,i[�b76��{Z�E6F�Q��,?GBs,3�a�������`���T�$%4i���2�M�����(�l)`��=���3���&��K ���3���J8��w��Aji�:H]x��D@��_*l���ĲN~����8= �r�]�l|p��"�|]&��Ƶ!{�����u�77Ya�wR.�0��F�H-�.P7M�Sa��2X�(!jF�nɮB�&u��]�E���AcA�J0��!��,����d2��Е΂-Z�>�d�[�an,2'ufj������A��h����	�"��5k!L����ncs֦<p�,K��iX��1�&�s���<�6��#�ݨ���u��:Ӻ=�p�2"�|���L���aBS��D��J��<�ӵ;�]Xd�GD��Z��
�9�c��=�_~FeƓ6 ��eT���l9�el�c�Pp7��&��S$�n�sg�Y­�XSP�UڮAe���[�lBH�k�&5yv�HИ��!�� O'p��#_8F�и�f��&�u}����B�*�QDQ�X%
��vۓm�]��R�
В�Ff��.Fѐi�-B������#�%�8Yé���KO1�{gf��L>���B����|/|���Ţ���CH�X���C[��q�zT�?��N�Ȟ�C�UK��g���0\4�N��u4�1���r�b;�{ ��B?/�ю& )H���e�Fi���I�g��;vE�a$%�����ܝ(�ݕz�I���Fba;�Y���M,G�^C���s�D��x�\�x?�d���?��O�8U(��(���n$N<�йA/���6�<����3��#�&�6~�Rڦ݉8���:Q�����柌��.�p�_�]�_m���W���=�t+ ^q#��Ԩ��#�IOJ]�GK,��)3.;D�r8["�m8E���z(Lĝ����Q��Q�'Ht`[�[��#%�AI���fa'�遀���q��e�+z�'�u?j+��m[�GRR�$������u��"��QMI/�mL4��x;��rU�k���*qx��GI_P
p���Q*���Ys��4���]i'x��h<9s�9����fa�%�*�8��4睿�#D�����	��@|��X�����~�L ���W��dN�����j8ƻG� W|R�Lz����j�u~D%�ȕL�(��$1��z�VNh�u��ʖ�˗�
��,���[��T�xg�Z�4b��	��m��.�vֹ_k1��tO�=���q�Hf��ǘ�uǅ;��Ǽ���X&n�X�r` ���̠D�X�6]�q���f|�R1�ӝ�麻�#��f��U�֠�L&�f\�}�!�5,�x�>P��dTd��S��;X~H�W��lV�QY��a$\g������b���&C�a��'�96������GV�[Mf�;���`+<��x�8ǹ�����7�'���rɧ�谙� �3�b4Yڬ��ђ�Y>Z�*�+_{F�瞊m|0y�DL�������JS����a�"�ۗ�	�mn��U�,})�Ϻ��L�����A ���j@/G�|�rˍo�u6�ѩ���rH_���g~�幋��R6K��`����λ|�.P�Ӭn��2d��h�C�1؏�7I���8��z8�N!�����8�@rq� �ذ��]�JM�!|��.ho,:����T%�ι����[�Hp�hg\.�3�ЯE�{R:#�bY\���~�9z��ju������0��|�5���cfR}7�	0Z�fF���V-��қ:U���m��I3֨56�|{ �F�(fh-	� ��{�>뭹�����Nr��J�I��Һ�o^��1��0��	��hх�3q��P��\�B��^�NmF��[WXK���BU�0--¥gL�UUA�5!�"|�U@��Y���Sg����J��|�6�o�Au���fWBQ������)����ӌt���)Հ]$V���O�����d��є&�"[t4f���8J�k&w,�d��STy�2ņ�\��?t� �@3	u�=^Z�aHMLc/8zk�� �>0���������r]��@��Gz}Nh(�ݧW��z�������z?X~	�C�~�(�}�R3����pV2� ��`}M��\8�ݢNL���j(ˆ�f7R��4����(UQ��y�P>�%��E���ĉ��7��~
��hr����%_X�w�"tƁ9���I���]Zȅ��o��3$�_�Ra4��Z9A�$b��s��|�dњ�0NAɌ��e�yH���q)1��m���EmW����8��l/E�s��2&�"���0�g���~.����*��UF�|�r'�{�bl���o��@�=K��u�E��i`����1[��$+��Q�|%��V|�������e@ЊU,����t؏���^��'�҂������[b�hE+;2)����c�$�Jt^q�4�ex�	��Q>u�^kJ���p� �"zaB^!o��x,*��"Z|a%�tl�����K$%�ZL3س�e<����7#|	�R/��^�7S���1vo<N� g�/�h���!�#ɘDh$6$�ցb{X��i��8a'X���槙Y�Xp�M^����6�gӭZٛ��v^�y}Xy����p�:�=J�B�>�JŶI����
(WK �_(��섢&-�K� 
�*|�s˗���8i��UKP���w�yH[r������b��8O,?ٹ�OO-�u���&,�,��vF�l���&Lr���_.!3�%�k��c�|M�G˾�`�B��2�d0��i��!s�<����I�\mDy�x'iT�7��EZw"�r੖=�����H�5�I'� ��3���"g�ݙ=kС�v��P�(��y��*C;ذ�A3�ja�PW��fQ�\[�h��U�ؘϳ�b�n�����{�P�:W���%�Wgg/tU�r�p�.v3q, >��Zʨ$��d7���$T�GI.�Ѳ� v���F�qN��
Y�z���r�E|w��p�w��?�-�#����1���?Q�'��,�r �uˑb�T#W��w�\���k}��Y������1r�1��);�[��r�I�dr;O\9 Ldsɰ}��Ln?��l�l�1eF�}�����p{����&�uv��)�e�sH�6@/	ы�JT�.�
"�(|К�G��ԇ�������ø��*ί��?��ENX��.�5�_�7�/�"暧w�tW�j�@e� !��S��Y��}9t*�<���pl��,��ǝΡ �|yC0�VB�&�����ŷ"�P8I��wf��2�	+[�I�.�u�yJ"����C��&e����"�&�7�»��b%Y��Z8��T%a8��d_!������;���~�!J�p�䙥O�[�P`�C�8U��v�J�pT�3��n����}���s�מ���`,f8�{�MS�: �_ll��.a��'D��<��H�<MaP��'>v��K#��M~ܒ��@�o2�건j?�)�Ck��Ί �jLc�}UyD��Ɩ�,o6٘,��'�ی �C��bP���д�x�9=?)WZlک����������-�1d9bw5|xF�CG����>�POnw����z3��c��<����?�Xro�&êgk���\{t�lT�#.
t��46N|(�e��JM|�۲eld	��-$������<���9Z������	B*
��jS翹[S+矹����N�M���ԊO=��s[o$#$U��?vgVf�ڐڦ[e*����u�Sռ���()�S�؟�R��Iw����q�������O��sWM]L#����
*���0v0�x^�\��$פ.Ż����[�� ;����q��x�^x���A��	|܃�s��$�������e��i%܆z���,d���H,��D�i�$�4��sgg��E21��g�x��A���,X���|C��Wz�~��&�檥	�4�Ѧ=�,�k�u[�պ��Z�F�wW�5�<��u�
���W���tO�U͜�e\A�6�4xM��y�T�l4Sh�5�A�=t�ߥ,��^�"d����<a�8�tq��&�&:0۸�*���(�2��M�#b/4�~���lu�aKB�g6�߬���\P<�̈́S6L�p���^qm_pt�H>f�e�̐��e���90z���J;�ǻ��$�<5��&g)P���˯]7�'��Õ�r����O��&�����{�-6�$��)�)K�ybH͸���k�*�~�9�]��1�S�]�pJ�@{������#!��#�yWd�P�w=p���g)�쯸��^,�VmlDR��|����-6M�����c����Co[����a�ڢ�SJ�溮܇~�r�
=���[���$uͱe�~
�C��v/ߕbp�;=�R:��&wt��R�@�u\a��(�x˾��dFy�1d��?��5�ቈ'O���&6��R����`J0����-��j�g�
��W׿�m�F���Bb�U:H�$`Z�?�t=F? �P� 2�H�Uj�(6W�Z����ލOUnh�3ìMXZ�l?Yʯ�!p@W��72��d��e��-���X����N��s��48��U\T��F���z��F�;x�b�v�M���
j�*�[�uOV�1>�K��#��SE(�璙&�WN)�ƣ����w�n
Sh ���YDO����Nf^����A�)Բ뫍�5Lv�Ƴ=����5��+��U$3jp���I\GP�L��/�;�2�i����SfV?�C�x����*��
m�҃<q�O��ޜp9?�9��cW-1�����Œ���f�?���rHM�S?�~�R�)Te�jж�c��x
�ҽ�ix���s�T@��|�?�+���P�M��<ΩJU'�A-w�{������w�WL�PgĴ4�(W���(�9,.#�R5GK�JĮ�K��9�iN���Pށ{�S��f%��y(1_=Nzo�g��\:t�>�_�ݏ/�����P�����	N>��-�w�����u{`���b�gZ�
X��Ґ����*�S���5����� [�g�G,� w�r����j
��GM'Z9	:�@�f\(��Z]"-�����ef&v�p�4��S�$~J{X:1ӥ=
X�����Pd%&n罋������>Zc��	�WqȑKy�p�+���1ǹ&T���Y�V�[�J}��]�y�I�%�宣�%�7��jg70�hzMk�$hOS=蚳�H"ƢQ�J�ʎ������AgZm`D���&s����bPڍn�@s���lk4m9 ����ʊ��{��\� �t���u�r�3�7��|��W��Лvx���|@���݊:��d�;�C��X�ϋ2*G5�F�j& �Sl�R��>������� �.ӄ��x���ʪ$�t켦�`���+�k1�e |�/䦋b��i�և�c�?��� �z�/��S3,���������e��i�G�H�3�
��].x|.M�Ԇ��.�L�xQ; ����2�p��ݵ�j,�gFu�g����E\���L�~��|>0��<^�ɸ� ��h�UB���D�$�nP��.���	��Tcbr�U��r�Y�#�e�z� ���WuP�_ɐ�:��~�l�	���PY����������[Ϲ �G̜�7�TI�⦷oʲ��u����2N���������ť��� /v׍0��{��a�{a�
�|lBu!ZJ؎��f��p^��ձ-�B�m��F��)� ^�_qx6f:>͊IV{�!E���p��
c}�A�@>Q���8�'~9'c��,v������9�� �H~b�f�� `��Q{��1���n]����5�A������-�KA܏��u *e��6j4l��A��Yk|�bf��B�*:�x[rY���OJ���P֭3)�T��0ڋ?��ΉU��A���D�5���4�2��^����v\R�]�A����	�z�}Ijx�k}w�Jذ��3��sHW��kaQ3�H����&$�
��u6;_�ר�2��v7k;�h�#WMO�����ݙ�j��d�Q�ǳ1JFZq*hF ��`1vXZ(���	��<�@��Ge�pF�|x�8W�V�I/k�ָ�I�B�vJO�i��@a+���?��]�ci,%n��Yp�=>��g���,��ԝ���d4�d���:7�/�X�����
�po�Ȱ��"Rњ�>	33�9���RPӧ#�g5�9���6W�xX;M�H�aI)/lz�7v� R�vd4W?��T �x\)�=�ޫE�,�H������e%��Kb�'5Ɇ�cnQ�mVz5ݿk�/&~Vߥ��Dw�^�Mq���6g㮮���X�*���]�O�yҴ�¤�Ygm�*HPo����	��O�(|X��YL�ISm���_�居'l�n@h�وs��N�-l��'�T#Sܨ�h��c',�#<뷗�}�����J�FK$�!J�N�sማ�%�Ъk�[j���~��doe�^�p�������t�&��]��z�<�Y���v�R���BYQV���c	��;W@?���� �ūa.���8.h��9j���٨��eN�3���.H[Ot�{ن��p�����H���V����n;2M=�_������ˁ6�[��k����!�gL�t4Z��D�% ��%�&�tژ��� v�P�M�_��;9����T���j����Sh֟1������l�6&��5y�u�;�P�3v�H����
s�N,~����Y�lT�H(�c>]J�ie^��N틛�sM�&�/�f� gf\���o�xC�͒��|�bHF�o��F2���|�r���,��������ѥ\ ��B!��k�MS��X�����$t崎��[)]?�ّ��Ͽ�1T3w[N@3��qK8�#t	a���+�*/e�2h�x���~#���(_}�zb�IʻQ�L�xxۺ1�E����g����ý����6.u���~RD4M����RYnh�xq�Dq����خ�\ϱW��3UWh��V�c+KxS��I",d�x�
.�D8���O�s_B����٘o/��$R>s�������d3��Q��#Pl�D�ʧ)gB�����7w�X��͈��CihmL�óch�T�'�ɯ�i�������G4�p����Kv��g� �����*D�_��oo�`g��S+
:�Ϝ���rГ��-�w�*1�/ v�~�� Fzǧ�������	��6~�,��<+eF�ܞM$=��wi:�ݲ!Î�¤%eU�W�7�ٙ���ox���y28��e�+�&�#��`�/�r�b�O�ā��P��#�7��7��oA�o������>��{2SD�K�J`�(ء��d�[��-��e^���\�G�|�"۠%'��I\�O�d��H��YB�$t�\�C&'��Ј��`��6	p�s�
��m��s��W^����y^$��H��g^Kʲ}��DU @����N
��Q��D�W3Lb�[n�dk#�s�7��S�u�fm�&X���ƕ�O�g"�k����'��8t��*�P�q7s�^*1k���Uaڹ�c�K�WuȂ�k&Z0�/0�����ٕ�A
�g8�*���(��1(h��P��5݀�mK/��b�,�������O�����rM���2�55Z�gȯ9���|������V�l
�����L}	;˞��ѐʴL��i�iҕ���	�������W<{p���;�W����6Nq��S���P��*'��`q:[j���-*�߳���D��f��ZA�B�|�K�'��m�Z�n��$�Id��=�I���r5%<��<��p�TǠ� ӂ�?%��銄5�	bB5l?��8�UNq����ؖXgX��Xv,<k0�\���H��i;}�E��y��֒Q�-��Չ`� $yn�l#���n�p�0��1��Y��}��)�)7.��{�gQ���ZK�{q���'_d�/�6[�6@8
@ �í�L4-1��rn3G�5��q������ �qI��{2����SN��,��P���^V�ހ�{-�H,[�!��o�`�������P���{���NV�y
xţd�K 8ݤ�Et��r�37)A������h��>j�{�%8�F�s!��U�E�q�>#�|���U��OWu����+r��\c�Z��q�3�[ӹ���KN=����/E:�ps�	r�Ç�"��d��=�%^�����!Z��ܝ� T��;�ÿ���A��ͭ�bw�����;����a������js��ī��*uZ�N;7��:-� H.�CF'EFˎ��A)%�5����Me�T��R��AȆ9���g���69d4+��HL�U�/��!�x�ևZ�,W/��N?�Zy��:�����r��yX@!�����(A��V����z+��o��<�t��{&$�WQ�dV�����I��2��3���^�7ؼ�q!�{�U�{<Oh\$�0Q7��:)�p�9��~t��>�w��,A�����9�j�5媃}U�dp֢6�xb؎�1M%Q�Li.:z����_�O��wJ�	�FyaihI��D����C��C�@�V
_��&S�^���&���K�A�W�N�$w:���#l��-��8�ajľ�JP��^�������Q�ON�$J���'�o�C��:DP=�_�H@���)��!'����������y )��<:��)ke���Ȫf\��&B�_K���؅�Zk�]�>^�x߼
�{ɿ�
��w����4TK#8��ą���2�/"C����#�5j�l^M�`��
퀃���QJ�\�ř�U�!�R�*��0�����1�)#?�_�F�5ɓ��fp����o�*4G �����?uJ�PN�ChnI|;2��BTre7yY	Xso�4�w�7���&0G��ŏ���o�sTGg2�LR����w�*����]:�#��O��X�p �:��r����1"hʫ�Hj�N;Q�X2(��/������ʼ� n�#!��T�rbUv��)��
��X��Z����xW�㠙�nIE�W�`�!�вi��m]j��0��<h���9=r�dYp��*�es���Ykct=��5/x"8�x�K̷�`=ֵ����)���}�Y���Vb��Z�WQ�Z(o S��T�6�u�dw:4��{���^n��ʡ|����C��2Hoٓ�� 8�;�Cl��
�랰4z��ݨ���"Hc%�^�g�~�Ktx��G/EQb�M���@��	^39�B��P�`"Z� �r����z `ENXO��˱}��i� "}5ӫ;��4I2����[�ų�#��?�Q�/�l!v�p'o̏L������쉕�� �9o���AL�63�������V	������Ɛ�*�:�������Ͽ{���п����:��]����}\��j@d����i�ۮ�5Mvc2Cj�j_�k�/�󢔗h<d����{.g�~��xF6 �������u��xU�H8N|</��%�x+�Nc������n�A��q"=��2��h(���[�ʭ�-���X�(9�˫�i3q0����s]�?D��+�=���?��L�23�U�_zcC �ˎ�������{��t�!q�J�V6Y�<��5��c�
oDQ���_!�wt�*���Q<^�Y���q0{v�a�:��ۍ;"5 =��w��x5$~�L��,�04�pz��.L�i�(B�ʛ���PG��0`�K������`�G�ֿ�F�C�	�\�*m���Im�'��^7���~_1tqJ	n���#rǫ��Y�B�d���R�8��o�C�"­b�K�� |JV�����_���z��E�[�~k���`�r����S֎���L�x�IJ]>l>@Fߡ���f�����y��_MYz}Qجquń�uC<P`���&P�"r2&=5п�����+��J�jCn��f�u�c�ȴ��l�0�H�� ,�T��%�lF�h�F�����ɤbjM�Lj���<��5��d�^�t��ʯl���~(���i��
h�]��-����@�,�ro�H��b�&���W�5bh|T�?��tl%�s���kv{{<������܏w8�<�74ޅ�T�-֏���=�ML׹\Z��RA�mgŅmcLwUg9�-�b������ !"mחƖ�Y�͹c.��m}t �n��ٰy�4�;�>+���C��#�y߱�;��E�Y5��F��$���ߨ����t�E��)km�V�j/>�P�ls����h�@��q����7��৻�2�_N�L!�\�M|w�sK�Rc���+y�;�' �����(+�0m���~��?�T�����a�gQ 3x�9�'Aʛ�*u8^�Jj��P�ĬpTZa$�8�AӖ�82�p�n��g~���Дۚ 85�ZC��׫��'2�m�?L�1��lʣi�I�Ky��--�
.�ku߽8�3{I�rEMD���IG�6/�����M���yAE�ی"#<_9AI���$��~�!>��靠�g%S��g4������V� 
ʚ��������Y��t4�u�K�7�A�(?�c�����u�fo@���(���@�r���ߴG�إ�j���
�3�du{N1Hw,�-0U��l��޹?�=
bv*����z������������u��|ڜ� m28m+�ɵ1��P��A�!|��ol�!	���9��걎U.8g���q�V1'�l}���hW�ڦu���eMu�P�>��lV����[�&5���[?�|
>V0nrY!�����^�S�uy���h=��8;֫�2�Dzhw��C�/�@�݌�#�t�+L-��w��,Y�?@�
lۈ)l�FI�ړd�f�Fbcb]]S��W�����9U΁�T��v���q��%�p?�^���;��5�}{���:4&�ۡ�C��
��i�ɳ�rU/�zv���o;��oy�T��e�7���7˸SiEzw�"�ԧ���YE
�ef,r��0Y������˒�����g)��r�ř�e�/��
F
F�|�]�9�u>�����,��0�$��G��j�N����=<���-���a��L��6���6nm�L?e����*�d������ �@#����(*5�}`��?+��h�FL���.�� 9'�贎2�سւv"���דE���|�c*��D06<羔%K
�6�d[=EW�FX��t#R�/C�`h�!���Uw���F�+�>��c�ժ=%�4�@�ζk��u6B�&b8Z���~$����Cq!ާ��1�������'����gF�F�g�ѣ	��:��LJ�����p��@c���Aq�Uc�+M�6ak�c������dE�u��
��evh+�����Y�z�L�.�}�A�.�hF��O��`�`ҧ�w��r�Ȝ3����Z�SI�st�$zOu�h���>�Z`I��W����H��ȯ���zM㎚����g��Ѻ��*> ~���f���j���2�[ ,b�i��j�B�ߖ�&Z�,���Ҹ9mdA_�qY���H���hT.�Uv�?����,�Lܬ-'[S=)�������`�;��ҩ+�	����h@[^�W0@����ӵ���r]�}��|��l�����*MM�
�	�n�d�d&z	g���r�ݛ�������X��$u�3D�U34�7���$����zd'�i07!>/-$�/b`�����tc�%�g��kD���6����T,��鍄�Χ�<C.2��/��@��g��8 .��_=����@��b��'�?}�-�����M=
��_�_S+�L ���k�P��Nx�R�C�E>4�\MD�$*���F���2|-}.�{u�/5t0�5�P���?]q�¹�����S���T���FÛ���<��K����ahgF�z+�p0��	Pw�,�k(�P/�	EI%q
8���֓��̱��c��|���ԂЃ���NiP�N�D���ȇ��C77�ӵȱ�Y�	?`�����8���)�涮>�g=��9����d�S��)Y�����+��_iCe5��]���p
�us���W���T��`�+���S2Ȯ���������Z�����8�R�;�\���@�`X����
�x�$۽�I��0H��aj�4�%�$�vd��j��֥%���(�
]�A+Q_5�oխ��%�i�-��A�n[ߛ��] �^�m�k�F�����Ş|л]3��O����CNIR=�#����]�I��8��r�l-�-�yT{��S��0|�9�R|KR�-pڙÕ��.�;�$Z���I�;��nh��Y%A�}�3aFi��Jc��>z?\#�|;��R�g8ˏ=�52�4�̈e=r��"uE�J�[���"M?�Ѳ#���q�Ɔ����E���SH�L��3����h�E��$�F �b����k)��0���~�����b���3g&���HӀ��M������W�p
��M�UV�^4?�W��5�u@E�̡n?9QF։.�9g{�s�Jum6�lT��������R�+S���l%�?���RK^b;��9]�̱�.%x��w����^9��o����"J���~�U�Z��k�P%D�v�jFcJ��@Q;��e�cOޗ����wjcNdp�C �$�F���Xz��4ޞ��.���񽐐P�K:Ӱ:�:D#�H�"��Tm����ɂ����lB��.䐈��QWCWb@��~�2m���^��ٳ��g��n7� 9��b���蝷��(��Ip2V���)���S<|fm[n��b��������ii�H�Eq�!���Xpz���$�>`su�yP�+:�����p{�X�6��U�>M D.���<�$R��iR�@�]��`]$8lv�����&t����c���۹aR������8�6��ɑ�2Oom ⮻��lo�*XA�iFO�4ϓl9�p�Ne����R/o�b��I�Z[rv����x�����lw�! ���{ǖ6R�fC:~�w�Y���~Sj���$b*����C��1�I��n��$�Ғg�I}��MW�D�,�E� �|ˢ)��1 ��uQl���Lhj���Ng�^�
�8y*��55`�I�Ll�D�W� <�O�\35z3�<�n� �������� �̿�c��,�G���7�C8��|[)�i�b��d�;G�B:H��9%��U���;�کt778����wf��>�Y��h��3�Vx��@A�0���3:�R���o�6B�77`�Qr�C��7l���?�#:Y��X��l�W0�1g�{(���<UF����qO��ͱ:5��~��D;
�a
й�0X�ɤ��nK��9P���B\�ܸ����[%��m�8v��C�i���Q��Z��W�A�~7N��� d�f*��&�%Q|�%p���ꈊ䞎���9�Iao2'U�Lq�ߍ�y�T3�4���q����"g���k͐�QAZ�K��cJ���|���L��{1��`����ϣ�u� �9i÷Կ���+�U?��qD&_��kr��C[�����x�)�`��L�É�5��Қ��^ ��cP�|�զ����T�Vi7��L�֟�r�;<�%6�	8o�f��|���h�hɄ�z���p����M~/��'D�q1�� U�JKW�%�5�/jS� ۹�/���Zg:�K#� ��D#G|��J�~����(O�X��L�����Ɏ�������ŭ��$s�ύ�gz�OΈ"��І�l�a+�=L���k�b|ص�Ai�l|�n\ż���W��Mӹ��ZO֦��\-=� U�i�=N�C߮�I=[��V�K�d��n/qȗ�tmQkf�(f.WR��:+�阿�hz���r�J�Ϯ�Toš ��3qM#��ƊN.��\������g6_�D�`��Fg{�n�#S�t@���E�q��w� Wͥ��a��2��d1��&��b�^ՒHeA���B;[1�F$yR�>J*�fQL1�^��P	��	#U�}E�r��=@V鬕A��#p�����&	�'��(�͚'��^��ٺFOٮ7�2I g�zZ(�̔��ąL�:M��++�+��)���^V0���|��>���Ȣ���.1�������n����=�O�J����s�`��)l^�7�._�`a{�iљv��k�+�-���荔��7�9ɹS��u}���m��"/�����>>������Q,�&����������d%���,���p�������s3��@�lH�m[C�Q��@�+�#�}���������E,����tD���ե�N�l0!Τ6��.��	M��Q�qa���fk��y�L��0�|��l5$�'j�V�"Gl���)���RN�z+Ľ,k������M'�M���r��~������5�֤^�������+��K�$<��1r�<�į�ߨ��暃P��h��OJFy�5A8[��	=�wZy�D�ץ��L��8�^.��Z��f#�96v����o�ϭ�$e�(���~W^F/���GQ`��?.CSh�Ɖ��azW/���]d��(�g������wT�a���H!a����AۃRR� d�U��0�{�A�m͌��'k�kC����R���W3k�g�.u���N@���Э�gNI�+"��8����wFl�b^�\<r���U�-�tT�8J.z㴨hź�����2��#,�Egg�gvZ{��]����,��<z�W����O��U���u�;:*S�i;�H��'�L�{8K�P�Z���9Uf�1~B��6{Z�N��{��`b(|QOM�q
���x���i|s�=]�pnD5��qx�k'"���Ag��x�^�aOp���ih��6r!xٮ?�u���i�����y�9��	b��(�C��gH��;F @ske�%$΢�|��x*{Y����0�_�pb?�?�Ok�')���ɗ@>=c����Jd4.�ͱ�I�#u������m����#��>n�*ό�<u���*�[�yE��>�֮�g�C	�-z8����Sm6rM�֢��"�k�zP�O�_��� ���5�b@��g������s�t�^{�t�?- �{��Kk!qiW�|^P��yYC��~��}���w[��R��!G�
k_"+,^��0���<f��u�M�����P�fZ���)w�}�z��&�����{�xc��Pl�~�	PD�{���bȝ:d5��ꚒG��l�������{R?'$���'�-=*����u51���S9V=u�.��]�G�z5���Y^Y����#Y�4���I�?G�$�ܣ��� l:���47 ���	,�|�e��?^f�	)أ�����V|�@�9�\��;>J��4ϰ�d.P(�Iӧly���=����%B!��ęE��M2�q��	L��F�W��R��t�\��)t��IU��e��y�ߢ����	A���ؿ4<i��!/��+�����W㕵� 5�B�L9�Fw��Z�Z�2��҉��|_�,���AGx4۠ch�cz~L�rF�V-��٥)�5�%ˍ���qsD@�7��r��b�$�Cf�Ik+�����<�K�J�Äz@�?B&%���eORh�3�c��Ԁ���~���0��ZEͰ`�E�J�ޘ���aQ��+ZZ�gRőj 2�16�_e��W+]窏2<v6��HO�Pb��CY{�)�7�j�ee�T_3�\�Oj�@�o���Z��i>�˰'d�W i��e�j,ذG^����V:Ͱ���f�@���Y[f	_Ń��^�np�;Q'dS.t�%�:����4��݁�c����Q01x�E�+�4-�b!,��Jݜ��ߛ5�dT���~3��v)�����*��4�dW����Yf?��(�B�^��Hy�k�p���9�Js�c����	�v4��l�$wz�����V:?o��u�ZXP��1��d^B�U����:K����s��mԛ��.��)ZM�D%C��R��3��]BgI7�<9L���v���gp��x2�?�E��҉k���f��[�A�L��ge������wl�-�?��rÿ��*83�/E7��B�~��.��LFʒ�)���٠��>&���o�����0���dBH�T�u���@}D�r����S<"9RF����Kz�ܺO���vh�x�I3Z�g/Fu�����P��y��N��eJ��{����B�����H΍L"a>B�?�-�u��Lj'��ـ"(O��w��4lW�`.UQ�"�A����V��}0����j+x������Ҩ�u�y}Λa�tH��~����zca���6�
���u�[h����{���ť�G_�����e^f�zZ5�9\f`�9��BO�P�9�
�R�Kw�:<��[�}����%ϧ�0�A;p-k�!0�=��Ri#��������i{6۲=�>�4�>nIt��bфR��P�!N�}��x�䑜v�:�~ͧ�0���x!E�$�ciG�7�F�(�_BF�-Oqwm�B_����᫪���ώ�l��T�*��O��@:P3$
Fs�����@���1�_�W���lٵ��6J��DB�z����6e|i�����:�u���輛h��d)���o�'���6������&��@�H�d�h���+�����Ul�T�u@I: "6]�;��Vu�%�h��w37x�qs��y��t��a�Z9X��STE	�A ���"�@uUəZ����S������ø���.z�%���ns�'�{���z�X8ġ�7�|����T9�"���B�"�`6����m��_L�|���l�}�<5�C'j�@������P,��rpf�Us�mi�w��<�M�^
M|���%������M���jC͚������>��-\�/��>Kp��Y_�,��~ӟ2�<��>�w�������#)z���H��7�3���m�a�G�7��Za��cj��]����D{�rO��H�!�wC�wuGMX]���c�;�f}{��R���vX�Uk�]�Pf/V��(h �~��'G�
��9��*���N�8��@�d_ы#�*�������ۗ�R���h�Cf�r!b���W:�s|����f���!^2��y�cp,�����w�̚�as�����p~<�.�-�^�̠���c�o�Y%�����3
ruǁ���+n|�+�O��*�J�`Ў~�O�(�"�>��Vvep�[L��q¤lDJ���7.�U�w'�(���0���9zcǳY��7}ܹI�������Rmvp�?lՄ�9,3,ݠq��8W/��S�}d0`��ȬE��*�b���i(_��\_[�D���u((��&��|߅��_�[B9�:f�z��@iX>�>bc�w��ʝ+1fơ������!D�	7+���!v�����Q����/cӦ��2��!���0�;}p@��e J*W�*���1�(���tR�)�>�ao4f7�â@��c�>��P"��:MY���*U��:��[�&���Ě�䉺�>h�AG�v�B�*Wb��j�b�t���l�U���)W���xf�O����ݤR�][35�ǖ�vW�i~ݟҿɠ�:���c�@�c����%F��7�	|�U���`�,����UC�~�O�)������6ׇ�y�=3��/��!�qcv=I�� c�����:�?�]o�q��m�Y!�H�Q�(n}����x.��+�e�q$�P`٩gnfs��kߡ�wF6`���RX0;g���C���#<<�k�VhЀyV�M	��dfGywV�����0��Y �
�� �G����:C��`pc����J�u�E_��J�t��%)Et�EMt	�)*�Q�js1l4�@N!6;2qs�	Fz�>q�䈎��%�_��@�uJ�<k���f�zo�fh�}'���؀?ʚ
��a݈y�=^����U��%p��;��
$�����¬�jt��tk�k.���2��z'X�:����pF�i�p���✼oP;p+{�$>CJp2��y�����x������b�m�Ӄ��N2?㛍��GO
��Ee�l
���'��y���S����c�nEG�pD��k� �9�7�rq,��SX��V��QU�X0�,搥�2�D����@z�Yƍ	���燭.�}�E������z�S�_C8&x)��cc�[{P){�ʤ��X���l��H�E��ѽo.
�|J����2�əmj|��Lz=s+�RC1�1}%���ݒߚ�_�8��{����d��?�����=�K�a7�66��Ȳ���#Q�y�\Ú)�!�����Z3w�''!F�q3�7�@�	T^�1�)˽V뉕m
_���H	~T�y�S�]�����2��S�0:��٭�vdV��4#��&�"=$�1�ܫ��[ٜ������&v�ȩ���̬��)y��Mԕ&�y80�L����C�0�,�t�ْ�%���ͪɖ��:��8[?'���fF�,C������AH�s����"��h����8$�X��\rZyblVR��#���Q���Z�rB�'�9��
󦳐����!W\���kI�A�^>e@�}_^�@_��J���%F�;5������4<����P�o�zX��A�۽s+���-0�\�%d�jMB�uV�_���pe�=�N�������`e��O�����M�Jgo����R�G�S%����Nv��uk��o�qNw�� B���M�>gq���H�H��uX�®Y!TB���G��- 見�2��V(��]�z�ĳ���te��p3n��2��~����s�>:��;M<_�ų_g��}3.��뵎�!��k��>^�>w���,wȐzʏ��+C���<�_C�4����Cn�'h=T��Pv�C�8�{r S��C��mڤ�E�N]\*�h:��+k耾w����nR�6�����j0�Nk@�v�PP�������B�M S��ͪQ>BR~K������>�uܾ,�.��%��/G��D���cZ�|L����z�jQc6>-���P � i�/z�Lޣ��O7����l~��lD�V�[Q2v��w���v��4� C�J�]9����m��m����L���x3C���2y��.M�V�'݃)o��S6N����z�����htg�xl�=�Iv]y9靪���*:�*��k�� ;{�A�0�B���lu�6�Y����}ᚃ@�T^��>�l>冖���8���2Dݍ?%�iȀ����T�L��m���A/s�vL�d��p�*f� b�fS��ˆ��D��wGY�J��m6�c�Y=���r{t��.�~-��L����#F9��K� �'U�/ë��|�BǎO뾙���*�5d��O�]�yg�p�NYK���u�44�'Τ�C%�B#�\�"Vi`ȁP��ï��u{5��&����{�Si-;6�"Y�A�޶�
�b��!k �1
��f��p�+y1A�&*��Z_���^����(e�ly65�������0D�Qc�L���f,�%Z>�iAP�Oʝ	��s�2�m����-��AکC��%`	a�e؞������!�,��ǩ�{pl����6�M��RH����)��8B�Yy�)�\�%����曀���^��LRۖ�Ve��9 �&�v�yX��|�����4j�o�pY����<��`�wR���?ɠ;��n=�m7s���^ E� �.���L+��B��E��uӻ�^��ը8=�� :g�\�y���(L+�u����4�k@3f-:�#mN�^ߏ��FB���h�z�ד1H��*�����*��0�'���w,�8 :�r��#
!�C=�}}�CA�,�+T���2�3d!�9f�S���QtJ0��8{۫=�,�K-���:��4�]PD鴏
��GτV��Z�Wї}�j[|N���n��,j�5^�9�P�<Җz�|�ai�J��$���Y1R��A��w��t��QY޿f�^�Ť`�ɤ�%�x-��f�>�����0UID��
.�+<0bOءjL��>B3���qDh���ʪ/(K�e>�QH����"GG����E/�Y�Z�}nmn�Y�q���VQd�����Ӓk��n� L>J�hw�?yj)�i�ڲtυ�Jn?��G�fU�E����}R�=y�-5�M*Qz(��oSz���������L9��F'o)���u/^�w�
�6tR�J��
e�Ϸ�����Y��#k�� c׬���,]�o�K2U�@O˙ٓyY;�~xL|�3�P��R����>���Eۜ���BK'��b�Y�7%2����ĲBx=���R1v[<W��z�F���mz;:�e.h���S�iX�ڐ#N��,�ǃ�V���t�T,+<�J��L*�������/��ߟ��aqO\	�)5&jG�d�lx����k�:����a��f�z���4�5>��}N�g`Ѵ�&�:&���G���i0�1 ��=8}��r@~J ��R��Q�#�4���6p�1z��&_Rد��HGu��
�;�P�8�`.g�i)Q�ěN.��(Ճ��!�LQ��_:�M��f������:%H�Z�M��$6�\� 5+U*�a�۫��5�{u��r0řEAU������O6x����-:����{͝����đUFj��:�mu��D�	h��Dbh7�z������O#�9Z�~����/����N˝� �hm_!��_��A���Y�z��(�����xA�2y7�c*po�SM��=C^ÂS]B�Ⱥ�'�J]�C��Q}��C�6�6�Z��c�r�/D �V _�J0	�U�)���iQ�^-_�߻��S{��%s��?��F� s�n�
՞����w��F�/Y�[2�ƚ���1+/{�i�_5b��������zZy���&!�������(�	|����w���zl[r�M'b`�Ƹ$_��{�Ա�ٹw6��Ѹ�z��<�����DS�(�P��\���I5�4�Kǟ@��HQ���t��^q�
rw�܂u�Hf���WE����]�6�hW2��*�rX5��g�s��tk�tE�Ue��~7N��g�or��%��%�1_��	�H���V�=�������p���@e/rȨ�'��}
\��b��W��)��<�
���1���JO�����V�fN���"�',�um���Zx�\sɂ~^Tn��������:̵�� 	􍍻Ě${U�@]"�%���zق͈Zp,Lد��l���j���ߞ�?����h	-]6윁[ݫL �r���i
eer��5�3������ܗ�`���.;��/e:�*7���|*�:D�<���,��#Pc&���
�{f2;;&���퀲��#71�(�hh�;"!V���9e�2�>/�U���%���_m|��J/&�����9�!Gt"v[{R��Y:��R�ȷ���%���}�5���nj5���!�	�k���Ϣx�(�*gt0A��6�8x�	����d��� �L�TܭC���+,L�����x�1��fZ m{l�o��8�{���::�.�c�"����)arO��*RU:��{c.�Y$| ��1�"�e�@Ls��5�k��4���6����_IQ�s�Ge�p#�S�-u��;��r��q�w�?r�Z?�!��ЮZW�����U��sX��������ea�w���0n�Ԙ��zo��tQ�T�M�cT�1��|��"Ky�A2KR0���{^S]nY8EB�;��H�Q�E�d�:�m!�)#e��OH��Pޣ��mtXkZ�>.��Ҥ ~���F�����$k�8\��mC���>�u	1M[*�����o)�s�ȏ�8�j$�61!��D{#0��� l� �'B���������9*BJ�7j����W.k�Z�\�ٖ6F3`�D��s[�6�vwIsHG�7��3l�Q����e��ר���p�נ� �s�37�xg�������B��)�W�Uv�"�}�a��C)8.��>�0e����7��Vx����#��a�)�s��>g���c$R8�⃒��%!���&O`<�Dlܼ�g&	�<*^��ş����4m�e�;s�꠩�\Q@��3�0-�61b�۩&ַr�n���l��qZ����B��a�M��&�*a�r�G�,.c}U��#�&c���l�{�ڭ�w�\kڲ���. l����+$��`���Q��z�1� ��Z���<挮��+w���hm�ࢩh8׊�d�����1ß�l�*��Ҁ�/8N2������t��=3u1�y�b�"����o�/z� �*s+��y����-�����e����	$�н#�OE�+�!@��������� ����'N���v�F��v�t�%g�
jg���_��T��C��V��MJ�ʢpr&��-��E[ȏ4r�&�N#�`Go���-N�ή��y����	d�n)����Āf�]�k\����xZUޖ�"�'�&S?H����&��C������.I�c�9�XK�;�GNb�+���K9b�D�j�o�:���|I,o�n������2�DA�Ċ%�^�n3��f[�<i��[jU��JTP}֕�i��|�����[��u��ů�6������:�r$�i��p] �3w]��;�:"�4j�Xp<����|5?Ӎ����K�ּH'��ws_	<jl����TО^���ي��.��5�� �k���$�Y=.�&) �Iչvd��Hŀ��)�穕�g�q�i��3�R��hs`�&]��6�*�MkD)��2�I��>j}/���k�_0�m(ݬ�6~Ѳ�GϏ⎅���O<�)
J0��DXߍ}�or~��a���}zS���4�!�Z�H?�%���+��<J��[�X����(;/�Ț+ЂQ�9���t��vd�x�[\��c���,�7.��W����H0\X�ڟGv�|�Y�Zo�[�A��@���s�@�}��Z�5˴�y&c�I��VT���L�c=j�anߕZ<y�FWܢ�qd^�ѹ�z�������ܭ��Ja@?�0�xđG�V)GM!N��5�����EaV�q��Ǩ?���A�E��qs�⿚��`���Z0�k:VC���n�4D4�?a���l��8�5�u�Ւ,{Tf�~�Ҙ��vp�ha/�� T�7QI���Mj/<��
]hQG��wY���O�E�ٱ���C����Xdk�p ��Ğ��٩����%.e�W
4���!����^��D;{��U��#�r\���� �sdM���̭����	9���5�3̐�;�/�a����R�~�ϊҿԇ�:Wk�͛J��^Bh�Z�(,f��z�mf��Ǭ6gvZ������-|̧ �G�`Zֳ��w�M������$�,6 k�kx��U�,��&B�	���~R��#�2s-�>�5�ƌ�L)vv�l��s�M�d�|�Fz���#���9� &4�?e�����<C)
�`�V�ؾ���ԯ��Xq�c�O?�O(1�
bE2�>��Z�g�ͽri�JP�g�!ƴ�Z}��\��[W�O�b/9)�_Vk8&�q��Ԓy�Ê3���-���t�D�Ϫ�h?C�]�_HT	f�&b8��U}=,���s�+�G��L���1|��Y��N�E���)�-<�M�<�m<\��.?(ܖ�\��Q�a�r'���o��V�h��P���F�������M�>��i2Q3�Fl���<�K��= Hk��w��5�B�O	�R�T�ket��&q\K�=�b29k	�.[�y��%4�!
q Y���������uR;�<P�\{?��j\�+��)v��u�S��[���k���~r����������@�`�7e�2�����w�kP8�޵�)�!��rY@�G0F�?y�qc��e�h�Hm=x���~wNb\�߈���ș�n3Q]47&p�����N,)c��y:�����/!{�(.i�����������ĨyV��.�Trc"�@LL�g�
euB�M�F�,�MG�HB;C�y��L����9�]i��O�/y	e�h���Z�<m�}y���s�VD�JR!�^�����܍ �SJk�Uj�׊����H'���8(	1�w�a����lC3
�;_��(Q �1������ju;Q��D"�vu�мr&�F�����%.�?|��`nk{*kh �dz1�3������3=o��S�m:CN2���$<�9�s����.�;g
�
Q�cL��z��*�B(¥I���1T ?0��pc��!���04�[�WY�K�f�ƹ����+���9)E[����㲷6��Cu�s<EZ��HN�kD�>X�yz��(��E����[��ɽ��􇗘/����Bb�m0H�rP�ǹ-xg��^Rs|��Ͻzs)� G����IsSGC�W����v���|@�kr�:Ӿ
2q�A�"yJ��l��y{����VN�����i���d.���"�9�B�&V�j��b�TofeY�A��&H>UZ�����8���؏�����^Pk���A{�&�*_!UM�nrf`0�����.���i�b�pF�=���|\�9��P/�� W�,.R�al�R+(+L��Bs���6�.L��g��oH���425��>:�9�Wv��p�6Ó�)M"���Y�4kd��A3�<�0�t�L��>O�P�h�)�G*_�#��ZC�l�ߨ�_�Jt���I��j��@"���k]|�f1�zC�~���'��J��dı���6
=C����z��93�P(�s�G�Z�Wv�D60X�HF$�Bb�ٮ���qv��EX��g���,��-�m��yM�Ѥ.���W����2�5o���b�I���������?���*������x���\�'�������.��j�nmܿ�!T���؈�Y��w�9ٍ��𘔸&[�<�j�_�<�n�߿&�Ǟ>m����F����|1���Cv�8}%(�m8��ݵ0W���#�Y�.�i�pN>��CN�o�U��������:�0�OTE\-Ƚ5p��$�Z�oP��Ri{�@�'�+	Ω�ۣ,2���o�Z�e������.�X�@�]�Y���b��f�W�[��MR���>��k9v3��/{�(5n.q��{#��X�T�U�U0���P- )&����Z�и�|���/P-������簲[�GB�[���o�ɼ���b�QM���ޣ�;��v�����R����M���h�؂L�Q�)�K�EҚq�q��-���"ye����_0Y�� �kE���B�^��c-������`UO�1��nxE&���H�9�$�{�������E�x#���F��yW'����<�{A�a�J�KE�,S��������^�������]͊3Ť9�C�����	�� ��Ts�U����	Vc��i״�Rh:t�	,�q_�gK�m����F}yET��>@���~��~���U������x ��U�:6���.�����S8��+5D"�]�c���c�RA�T]���:/&�d���H=hp��O���ꜟ� �n�a��|�۪Fw�-��^��f2H�.��\<kV��f+M��ɦ�zGXqK> � �ܚ���+�Ly�B����e�44d.2�Z:jMm��0?]?A��(����0����R�utzd��}DML�
�u����LLf��bJ��.�6���-_��[va6A��O�v{w5:�V=֩��m��g=��Cnn;y��eɐ��<�N�sC;M38�=�Ä�(�����\	��q}D�S}����  E�!���1Y��`+�gZ �Q�.m�n'��pL�.L')?kps�} H�Kn��\n����JM�~h_�c�lk ���1>�4�Am��٬*-��/��G�@I(1}wZd��x&Lrq"�\��y�=uF��^4ҿ�:�p�R-#����c�I3�$��1�Smz��x���8dԷ�[�N��GdC.�_ ��&�S}��}8��R�!fN��}My=�u���;��7��j��c����j-|E"y�\��j�������DӁ��);޶.Մ�h� ��o��η5�����(}zHt�IR�����U�Y�R4П������z��t�ܧO�O��+a�ʞ��k�!M���Ŵ��p�̡0=\6�]�!n�V36U$�.7ds�Mi����O�UB��w��b�:H��,��ٳ����7ע�y��1C5���޺'��5J�v����T�"���ބ��*g�H�2�J�n�ƍ�R ���OP��/z|	s~��Q���'��v�3�ώ4�=�-X���i��:�}�x3?`� 5�?`Y!�*�J(Q�Hh����x=�H�&�>��Z�j��|�hk�zv����433�2��) ;��r|�"Np�rE�k$�'�N�p�� .Uc��ג"\���4-d��`"V�'������}��dJ���Z���ZRj��*8J� ڥK�<㑃�zxh<�z��1gȅ>'=v�]��[FCV$6W8G0{�DV�؃��T:�`Ƣ-R��4='�����uS{ט����%\#Cq���T1��襌��u`W,ё=�&{së�t����b��F�u���r���!��Y��{0d���8�~
7����8^j�BmP��A�i�Ȕ'�;<e�R5���LnI���Rv�,S�&%�{I+Bb)K�T��Řk��a���q�_~>���_{�Q	^S?� �N�b盛��Z@mkt�S7�ʄ�t04��M
��Pa Z��/}�ޜ+��C�)f���77E��Y���������!5#eg����4'�om���Oqُ������f����2A��4C��a=�.��#.�os����� /�I:H�s!�$�j���z��ʥ��@�~Y�7��O:V|h�ż�����R�o*���P����PϿXM=m��ʺ=�ͯ+ň�\eW��K�A���_�����WJ�0A<U�"~a�>�)33�ÿ0�x�U�ix�5G?l_��AQ���Ӳ�s����WZ��wE��� �z�-l�kT��(��� D��}�إjkW�[&�n�6H�������}n�F�
m�֞!~3�A1�����R���f�/B�P����8�Z� 5_�l43Ĕ�^�����_^�f�Ξ���uLڃ�/�EP4-�)�H&��sg��O�3-M�?��9%H�-F�ƆᛑaBm�4��:�X�M��ߏwB�_}��?v��ze���C>��{!�=����#�d�c�w�ǇK3���M�/Y6��X�.��I��5t�r��J�d� W�j�>SE�0����Ŷ
�H�@��w��?TK��c*UP�5e�/^���� ���Մ2Y;�ex�l��ٞ�$t8����W�?ދ�+�e���am��*/ٽ(�p4l��;�ρ���E�Djm����̫���j��(}�@9'�ÃAг���o�?39�^��Ky��9��C�P+�$k(7�y�u��ϝ��ez��M͗>iH�Xh��d�}0��ca"��) �N��l��;�:�tT} 3����-�+3ɖS��5�f�z���O��`�������I>s�i�V���w�OZ�f$�2��@\<�:��K��i$�>G�m� D-�50Os�=���ƌ�M>�֊�������wHR��Ϯ=����qT�/Y0���a�)�WAX �U6
h>����^�;R)�5�6y�md�}`�v�2v�}�k��9!�p�p@R���|i��V�Zs��VwA�()���E��cjMB@/q����T��{�5���Gy���5�`@�3Ⱦ���FVs�~����/��j�G�z���1im|�/��1���GK�^�e���jׂB����-\!
��YK�g���L�f�i��mG�����y��Ȁ@���2P-Y�3���"�!��0��d;�|om8��
�D�<�w_����F똏-m�M�)��ĎU�I��D}�TE!9dS��q7�޸����0��_H(ٞ��U���ǩh��ʌp��g��	PMN�R�Й�٧���?�X��n���1���1��#UH����u_{+���s�^�2Ј���9����3Ӵ�x�(ܐ":��w]\�I#��/��8+�}cWj�s��Y�e���<�Ξ{�A��p+I�Ǧ8�bk�$��<%Z���	�viA��}�m�a�V��g��^m�76CLl��Y~MQ��-4����ww]�FA���pIo��wTn2}.��8b%#�<.b����s	��J���J���r( \���0�j�W������Re�f���ۍCl�E��v�U��dp�	��<�$�tT�������,��&���FA1�l��EJ�t�y�"6��0�@�����s���e ���5"���ǏoCĭ:��7ѩ�jv��L"1�)��`��8ى'�K�)3^W�s'6Vi��~�F�M�H
m��5���݅�o�A�Uy3�I,��B�Ap��bhr�Q�_e���h�;���P(�N*om��~�a��|fN�%�&���+�r�Sc���y���x���C������F�@��ڽ��~����`S���"��
P�Ø~ac�fa�g��>p�1��Cu@���6��T�V�b&��j7��,,UV��!����:�¥��M�q�I��(ꭨ���ǰ���
"QF�F�|!����q)����:.6��hV��x�}Si2"�Z��zu���ZDo!R�q�s�J_Xu~Q��e�օM�;9�����W�qΘ��V)!��Քx���~9��0�y����H>lG,^�ΩeZ�Ȥ�]bXgV�5�l��Y;�}�T�£e���E-P�ϓ����6�R�p�A��F����La���3j��:��r�uB�Ԥʴ@YTWXd>���ɼ[���a��~|�SWc��:�5��!���
���Z��W��CJ Չy~^Sr�©�	�,t�aK���"��zLt�f�CB� 3v��T]�X54\LllMv�-��"Z��?(F$�4��t��= w�j��7��XE���	O�jQ�; �ЉO �����̼�/8�jnl,� $k ��c�_�N��Nd����cm�0('�ZT�~=uV�ݨ��?O�*�81�f��$��[��d�ؘ"�`�Ր\4|T$։ /�q�˫�
 �SB�<_۫��A�[���|�h{l��k�^&���EQw���N��f�F�;�+�`�M撣�v�������L������8m�*��d��u�kk�n�|(ý}C[����px>\����	pK?�6{����.��	����ƣ�f2�g��Xl�i��NfA�M��N<�0��L�[vV�����.���l��C��#"N����wЙ��ON�g�\�����	�Es��!�U �Vh�~ p��{j70�RTx����"$E->{@�d�rQ޵�'R��@�i�~���k���U
��y���?>*�k�\ަ�EZ7�"} �����M�u���u�6��?T����Fɧ �}k���c����~$IM�����~�刨���@���~4��[�&�`TI0� /'L!:y����t�-׀8��C'�	�\(��S������;}�q^06���gQt�X5�o�Um�$��7�!�J�D����k��Hi���>��43<�, ӵ ���ф�����K#��߆|�+�=R��߈�Ա����0�I���{\3��A�Q^�y�Gu	�V�Bkr���U6"�<�Fn?���X95���Y�N�M��O�'i�_Y;�ۑ�W�#������8K���x�]a�t�܆?fJ>ğY��;��+Pm>��ip �H���7*�v���@� ��Ɏ�t#I���o%H��dNN��u8�Mĕ�a� ��H�A�����	=3$��l�>�aYc��l��F�g���QhǍ|����crW�hr�/\��1����e�^���]H<�׫����_��L��-k�ɩd�A]�7�^� <����J��X����닪E��W1m��c����$&�ϭY�F#�sYea�1n5(������m�����~)[��`y�HC�^J�=U\#���H�.�h�Yй�8�J��pɷN@�gBm��-B�q^���*N_�lC��c�_�(��k隨��9hIm���T��^�� l�A�(`��%/�la��:b�5��Gm
`��#9��e�8B�ʁYu;�f�ׂ7ð��\����g<g=_@I�dv2M�&[@$9���$���u��7��~��Y�^E�g��	��w���x�A���6��9�33�u��� �)���i�5o:-S�[��s1��ɣ#��j�������f[҂b��}��"�KZq��((f%4E�P����!���ѭ�Y7���eG`a�;YI\Wٍ ��E���f�o�e���'�ʗ�$+lg8�W����I:��Ɣ�'���q��Q)}��_-��fWs������X2\KZ ������1��@r��0n�r�%
�1��#	��;�>�_�hm���/���p"DZB�p��|���'|��2��
��+��+s����^R�x0�cC�.�gR�GlT�{h����鼒�E�"��B�`�u�kZ�|�q�K4Mm\g՛�?�I�5��	��B��O,����HK��_&���*����L�0'��Vif���D�i��.�L�_�q�Y�"ڰ��#�!�J����pbqIA$o�7��U7�
�?����˩}=����qb}���2[���ǎv	Ј�o�[��K����H�X�iMki#�xX�:L弁}�m��?�tZt�\��E�t���AJYԈ�J�BhG��O�r,j��,�Qii*��:v�~�8��{iD�	$s]�GQ����d�e��ȓK?mx㦉8�f�F�E0�/積�x=�8���RC�g��:�'��C�g�i�9�,l�y�+(��	燬��i'�H3;?Qܗp��2��6"��ח�j#���.��"#��h�ӕF͎hCh��ˣ��
�/ "B=��I����q���)Ο��̻I�e6:덕���,��~�L���H��4v�b�!�y����d�}���ǡ�Ƶ(�B.�u~s�ZCk��,1Ĝ2�Y�8/�w(~3�n�e��7�M����İ�p/�	�d�W@]]R�i)>�%���푚��gJ����^�\��w~����* Y�W*�~��~ߜ7���!�Hy�b;��~�L�ٍO�J�\�=[�v.�`�cû�����"��ni��?�23b�[�]�=t!1Ô�����7�z5���,� �_�"FJ��q��>6�<�m7��ټ�*���|�r��������	a:�(j���|6�ǘ����HX0��P��MN&�e�8�(���ݝ!�5d�(6g c+��g& �f�l�b�هB�Q(?즏��eU�=�\I�g��!�0w��yfg�lT$d���M{�á���,����y՛,���r�m^�]���<mU���b>xBM�L5���x[Y��������o�$���B���AG{��!�Vڳ��ȼ��h����)]���sl��$�1�>G���&ǡ�Q9p�D��2d%�6����*9<��s���	ZMlh�3r1�;��p�*G?�肳
�xH�c��F}���d������!8�_��,����)��#��^���Uuh&4��Hq�k�Fy@
�6�����1;�p!H����ú�6�A���n�ӣ�r9�XZ�x8JG.6f�_~�'����0����&p��lj�����<).��4t	Q���x���@Ieg{m	��A���t�Hy%���4��B	�>�e��N� q�`�1<�Y�Jqi��vԎ���ȋ}��I`�}������Γ	U�}+�^�� �FN�UG�����s���9�|Kf���d48ڑb����˧'��!��UmE��jG�l�=ȑ��C�����G��۰��v���L�
y� ��
����\�N�������}�,�1�=wڜA�s���b�<��EXSk��P�Z���R��Wq)ˀs:Kl��M���p���n�z��ɬ1DX©p�ߎ�u�[��|{�|e��)Ql������SL�f�f�j�P��y� *����c(%a�qz��\��Qv9�Yԭb�.O�B�/:o5j����ze�z+]��)٭>~�<�4OЫC 8{�Yư}��ߗ����	t��&�j�ְ��N	��T�BG��lK���B^(ǻb�Ȉ�_$���-[Q���t{�g�&�H��R�3��2��	��.�Xę�\��J�7K1^��������q��]�.����iJ�)�]X�<�{�����]���)8y�V?��3�(��=�NED�S����a*U�!���l�b�?)�p�Qb�@Q�!�D�����\�����Q���BTI��4���'L}���e X�����
U�;���6F��:��Y!�T1��`�R��=Rj�5u}-����]��ݽ=�d9�L�ȶWlO���l~��	e�G�1�$� %~I������>���z�̵�	'i��m����Y��E�՚ƻG�]���Sp�� � ��[!`�(�Jj0���$��2xg��MF i�v����ݨt jن� }{��zKTɉ����j�L�0Hd��� ��P�
ԗ\��Oq�iو���Dq�$)�0e��4�P9��@$�DX?��~��� ] ��)�칗�9�>䃎ǧ�j`��ʌ�'0�ϰ �^4�g��_ѧ�2T7o6�Hh\�&䩏٣G��4��6����FD�U��[���_�|���v����W�ގ��)��/��v�r��$h���jĆ�˒�?�E��"�ʌ��/m�v��O;�R�G��f��O�$�?!Ateh���d��@g�z�D�X�:'����i{ζ��@�`XF�,�?�ٯ��+�Ӭ�Gq���l�h%��e���fS�5�I`��=�0����T )_�{���4��j
\�p��<���aW�������r����穜#1�V_�V1Q�2{�%�O;�՘|fJ<�K�������B�0����
�z�2�J�k��z5%�3��M�C��^b�q�QG����C��~Z.����x��,Y ���f�\��l�V��;�O��4�sQ��m�Z��>�r�E��Bu)��!��AN�w<�X��7��Pe�۟�HZlh����7E񵚦�B�ZD{��G��a��z�,�K�j����Ż�CzȾ��Iy�TԣXI�\\?��svߪ�+l�]�0"�˹��Ӷ_ĮԌ�*�pA����qr+�6��)"I.��m��A�����IΏ���5Nl�?M�:S0�c�#��P�蚣���
L����ڪU�K��I|>֬Y��#9�z�Y����d��Ѕ�+	Q�ޚ��Ruq�k��+�9�Ũ(mɋ�[�g� �)���9YW�OX����Bl�Z 
u�8I��8�G��+_�U�s��tW`�`̩RI�dlHH#h+0:�p�"�7a�Ԙ�\ݗ�dL�	�f��v�KT��0\�A�����4SֆDAc;�s�$��>�D�[v�9r�[�
��3I�'Z"���y(�h)��m���Ē�c��S�B�VȫɈ�%O�K��(�o���4.y��߷�pPt�J+��*AK��CD�rIV��A:�rT��xU��b�۵=��ë���"�A[7�>�k�@Ӥ$���OCJ�w��P�ZȟU�T7^�I����_���$��C���nں��'GI�=vF��{������5G���r��.�ǿu�t�����	�1� GV����4�DϽH]�gv^t說����)�| '@��m�����E�C��f_�\݃�~�Go�@�ǒ�g.2%�#h,d9�;�v�f} 0�V4������F��+�ۮs��lpEɿ�=�X�c��C�7TF,��U�i��a��)]7R(��]u���y���>���>�vYXN����MhZ�N�z�E��pMDz�._�>B}�,�c	�h�"'�o�^�-���J��W��k�R%��@��G�}����n�,�:_E,�~-��QM@���7JK,[08�l*��O�t�I����/�rC؅��c��$k#�Թq��9��`n��$�{��M�p�S���z>J/s#�ŽDD���c�]K�w����`���|-D�VW��[��A�3ȸ[l�+>�.����Rsq�׫"�cn>�B3�y�U��=e%d���*f�P�HxcjN��_]zS�z]d�>���U�c4�#[��礅(���	6�t��V='��2��A�Nϳ&�A}�l(�=u��� �[/9^d$���{�yƠ����	Il�T̈́��ZjC>�v�򒢫 ˵�x��8<HM��\��A��bh_�����ZeGĈ:���!$t� �*N5�t��"�af����Ɉ��w-��,VI Mpr	�@�p��D�ڻ3�cfM�-�
Z�V�G�	vG!'B@��8��]�fhL�\һ~ֱ�ƾf�v�����zA�.�W���'W^(ɨU��!W������|h�6/ߘI�9��Ƃ+Z�y�ą�!�#$-�Q���eo�*���f�Ҷ��������w׏X s��@h]��ǳ����/'��ק�xૌ�3ւ���� ��{iq�{�z���k�1��C�_*y���UFڶG�	��=�{׆�q��^K��y�f�6��o�4RBN����c�³Dկ�71�/��i���K��<� ����R�$���4��x=�P3!��H�O���S�D���~����O~&���a�*�(b�diSO\��D��𻮨wI�G6B*Q�4Dы:&������g��B~���ogUE�`2�r�W=�$_��O:����o���ͥ��;j1��}	O5?M!cn�G;E�7���v�S���ط���9��"Ʊ�ؽh(�J��b�Ш�)-�XTJ|�W�ܐ��&�i�|�"�ҷh�G���̛���D(Z�	��(��^��1�$�Jy�t�ť��e��v�����[�GywE��
��
0h'�~!����W�G�p:wfR��@	��J����d�j�IZ�Z@η���`s�������@�.�~���e���YZx�t/����#����o�Ld��l���ĉ��
n�]Q�m�*}_���Y�pe
m���_Ǿw�7}���1�.ېa���y���~h�	A.�����!̘�0%����D6�� �6���'0�n�m��*6��b<�����{�j��
`��:�2�H9{��Ն���y\6~1��t'�	&z��m�:O���qv���(�ȏH����Xɢ��2��]��.���޸v���~Ģ��;K4�����X �'?#����[���B�3�Y\�9��8+� �0�I��n�T��L�g$q�Sp=�9uYFqk��^Hd��'?Z(tv�/����(9ts�X�0qR��V�g0��N yǋ�
�r���f��ni4����U"\S�RȰj&ܯ��H�p��_����S��Qi��Ad\�N����>C%� ���iWD�X�`�E�66pů�N��l�	�L=� C���*bC}�@R�!*1����a[z�#�/9��(c�O�N4A�������@S��qQ��Pқ���
��+N"��PGN�>I�)n&�ދĬNDVY�YRK�t{��6��8!"������k�Q�����Sz��Z`&A'�JF�MАe��|�������.�~�Yի7�d+�Ҫ�K�U�H����.�����߽44kb�5GӿÏ}��yڌ�m*����4�=f��5����{�H�";K���YK��-�<�+��)��|�!X�)���}�`���]@����E�����kǙ��1�J���5�����aH7���=�s�;4G��B;�z��A�
��u��fh�}�����Mǥrk~VT��<�|����Iǲ�(�fY�R������;.ۻD��ǒl2��
�K�OuDVV����
]�*��װ��s+cۉU\K�j�Q��Oj�~��.?rI�~2�v=D�@����<��l�ضZY{�S�V��!���VJc�
1���!�Qo&83�b�f��VW('uXj�wz�O7���Q(7��S�LjR2�$��4�n�m���\��]��p��K�D*�(�枑s�p�M���R�z/�l�	1��a�$��l��by\�.��c���ש��Z`����f�L�6�d
��s��:�䪑X����H�ڴ��S��.�*]��`�y��6��Hɻ�;C欿�'�UR'�����o��
߽�b��H�UwK��}}��J�~���Â��_4Q�hOԲ��;�t�b�N �B��(�}���}�+��q�b��& _��ڗ���M�lqe��uʁT/�c��x�I��)�a���[���A�?!Z�B�F��0y��0D�At[ܣ>�i�8��6С���o�}���MV2)I^\������"�T$8�P�(��52��B��\K���jq�h>n~AN�C&s��myM�)�V򷼸D�f�>�?��m{uC�b�K?��Z>q��������g��P}K�`��b-uWv����Ti�v�df����t�p�F�M��u#�CY���:~�M�1�R�"m�U381���y���C����B�ث$����v�����m�9�����l�ަgQ��o�c��A'.�v�]"5Wv�dx��R_�T� �xF�\|?>�<Vk��lB'&�	�n�]�n;VV�2/�k�@=���4�r32+E���q脻��u+y�mg��?���W$720��K�MT�Ę�2e-�x�]�E{�������A��K�ɴ��D}l�+�j9c� D�Ǌ3y������Պ�������*&�W�4pJ���8F9 ��)/w&�]��If�)߈��|:�8�j�E��%�C%�:��Xe)\}d/�u���XU#�6�
�
�a�3��q�/��%J��-"͇-��@��"���һ�O?"���h�8,���f@��%[��1�&q��j��H��+
�&[M͈V�)K|Ѵ�┉�#��ov,���aS���lڥe���@���}0; ���Z�k
�a�Z��X��ͥ�F���iN8����7T�ܰ��]�7	��PBL���,�c�p7K}�%.s#YՈmњb8+�U^*��
�x�۸#Z��vM��Ѩ/�������W$fH����6A�n�v��w@ϔ%��ځGk���Wr���Ӽ'��F�I7a�C�B��Å�G�^�C.6enյ��y;��n>(/OՓU*f���Y5xLZ�e�<�i`,�|`,&,p�#3u�C�:���	� �w-�u���8��4�~'�͖��^W�=�A|� ;�{�aKh�u�.�cs�k�cxz�$������<Eӯ|��^JSΟ�����+�,'�V�����N�F���;J�V�^�o��/�3 �"���XqƩ�Rl��~����0��C_RC�G2x�����i����0�q�����MtÓ�	'�?�@�c\_���w�Ҁ�zQ`�h�urs?��(��ԯO7��D���=Ė}.� &-�Y������=x藣�t�T�;(j�ي1,o�Z!� �8�~�[�B)f��-l�X 3�6=I���\L>�3�~��uyy����ԚΚ����8i�8���ꭋ�0N)h�:�\^�BHZ�>mW8��� ��#�~}��rB[d���]�����յ\i|�~�=�Z�J-+-���ԌN|�LvM�ui���R�:����|_���V���.�ƿ��ζ��z��r��n�i���|r4����Y��"d�C�柕044Y��X	�H��pM���1���?���b�V��Z��X0R8^ ������{���pT�X'yo �T�Ȟ�CA�m�a|��~ �~b���7��VNd���e�Cd�:@[��c4�?^��s�ڇfmmy�i�xnB�$&��w� ��k�b�=	-����X� w�!��9�#B��qsx�f�y)M9� )>>����~�_�|^�Db �k�� ږ�C	�ӗ�-�<�$�D�������n�AI)M^�gY�4Η(W�M $��榦���+k����P�J�e
�QC�-+	�3�����*J��(��n�z=�/���՚�\9�����->7�Q��Y[�`�٘�h��ز�.]u��:���
�Ueü���m*�"=wm|*�;���{�β܈��h��:���u����\�2�&:��;i3�d�{{��^*L�0M��V���ɽ�	;���^xY��h�R:�i�_���b�h��1���U')�W�Ŝ�s�yb��d_%����T�� �5���F�������=Y)T!���z?�a3�B�=�U��OeZX��o��~��$�z�.'K���k��0>�%<�O����B���n�)[�(~q��Q<`�I,�A�����x���V���/<�'|;�����q
3O�}�]�3���&��щ���&h,���`���;ǌE�4$����pWS���v����w?��^��fQ���Cͳ1'KS|�ד�RO��o9����)K�3����"]J5�Q5�V۬0(h��!�cw�`�4�U�D]�>io3Kk���Z�^xl���+nV{�"���ė��q���U�
�os�a �TK- r\1�%r�]�y�w�F�L�,���L�w�&`.e���.=�x�Q��ƕb�{�zj4��d�k��܂���"D�92��l��"!�Q{UPv V��Ɵ�.&q�`��i�<#Wʠ�I-�@�"�B�5[��[���K�?�~z��ga�)R;�_O���V�q�����KW�+Qf}؆^�5����l*1%K����J���)��',Eq������TÌQe�{�kkP�	'�� X7��a�,��wj���Y:�C��P(�
E=�5��Rc�Ӫ)���~p_1I�u!��j(Q�������q�,r���lR�g+κ��i(�>�_�& _�)_(.ʣ���.��eM�F'��K/�=CVr+����i�E��0�(����0
�Ƙy5�vV�Jg͎���v jA�t��Y��+�����u&��""�������k�00}�=#��(mHc/�R�#�T��4��;,ѻ�7�����p�<
�#8Pg�&[��]#��=䅰�p	�*5z`�n���u�\����M���"������
�����c)�T���[��	�X�-�rĚM��#Ì�/�8��� ���3��QUM1b��0�ݤ���	�}V��k1��)��x��e�&uЭ��>ґ�|7�(c�����J:��p�v���Q}k Q���'�oq�A���
p�� �:��h�*m��ЖJ�`�2R6l��Z�:��s��q�#�E, s��Аpo��XX�4������N�K>�`@N������M�'��j�_�-�'�����h������*k�5��"�K�qWD_�X���(V�T��C�u�������G_0f�_$4?����N�
�0����Y�s0�N��\7~��x�b����F7�j�����{&<E�q�)_�b��� 1��/�6��z��ߩg�&�E�m#F��I0��%��!�Jiڇ~��s"�s>F��(��W��@%�B�!����S��F 0�g�š�s͉Aٕ�Y���1K�L<�M�Wr��B���(��G1&�/mn���$�����z���{�d&��	c��U���]_���C�z�-�2ڜ{>R�4��P�F�l�)�Q���L#ur"�d�%@�o�\R�k���a�x�'�h��ݘ�ʜ���MjG������*k��$�L�()��'8��&�;��/|ZZ	wdn���ߢ�=@���:q],P�ڍVuB���g�R������g`(i�kE�=d��\K�>�G�7eN�'*B8IrE��c���iv��;CI��扚�Yw�'�v����Hg���nǹ��}�_y۝%���"�/(6����ce���d�!��!�sU�/ꐁ[\���R�F��C�C�KH�R��8t�4�Z6{�wD��nؼ�4�Agb�Θd��qhU��}8�ݐ�}]�:�@�%<\�G2��[>c���P�Zl��F(ڑ9�Ĕ�������d�	���[���P"��	�,�h��SM߉�(!:�{��qN��wLi��͂������[���.�4i��&@��No��g���hR��H7`��)/]ɵ���H'U9�������x�&q�m^�Y��em�w�^���OVmq���A)�JH�'o�E`�������͖��q�ofvȴ�qʹ_R����
 }��2�1x��P}%-������e��S>�Q�� "�,�����l���9%���-�{A_�j�e�'6�RV|^M,b��X5
����ɯ�G��0`��|�JN
����\���H�>RƸ{7'g��q�Z�{>�������_DG?�V�G
B������bY5�~� h���|MO���爲�O���{#X�F��m.��d�l�����+B���H9Q��h	�ۤ��a�@(.n?���/�b��ˏT�x�b��焢1�����m.+�%ׯ�C����D��ϳLD���넉Y��ك2���zN$�Sc��ej��XL����9C�Z` ���c�vG��.,쐦����*����l	e�&ß�gJ�C�<�J��<���Bwda��_�&?�6�<�D��AK mJ�G+��&�c��� ^ͨ]ݴ�%j���.s,)������xH��?m	#� m����S�rq����lsg^}���ʐ�a�f_��>�f��=����3f�}��`�-2��a��^�d0�s2���gZ�l�#��Dw%�e�,���`�1���X�0�\39C�]���v�ԗc#�Cn��,���]b���L^��Ö��=��iv���U��S� \Ɍ|�}�������B��r��{3����hme��ӥ �����◛����Z<��UN���5:�|���0�ů3�������:��$��m�W�y��y��`Yl�(HL	#`ij�!'���""�4�;�ȝ�?�# ���%m9�u���QF��G�+S7o$!4����[����ܱ	��3���It���Y�FЛP:zhZ�� *��J��-5�&�b�1��o�u�n�<�Q3�T���"k|��k�w�d�1�$[~sH�k�-���\Io%�wk�s�]Lx�;�{�[	�hp�j¢�"??*x)��5)"�0�ǝb�Yg_y�Y�"��?���{�D �@�u���M{+����3(r�І3��Y� �����'�Z��5�י�#��k�ܿ���D��6h�Ѽ/�Sz�cu���}x�7|*k�(�,n����Ncgç��Ys�Eћ1���g8J�
Q�\C�y�Z��[wěbx�Fw�Zv�G������t���dt�&Ry	�j�F	��E��ط���S{!�	֍p9�H� x>�?RB{}G�%.�g�\3��F�A�'��C���4��	;zeTN�/�2[uG���~��X��)2�PHq��lJ��j�R�؅N�c-�������K�L-�Us�H�+�j���c�MĭW�,��r�y�?P��Y�CC�;�uO����Z���k����4Tә4M~T�V�4���\�d/����$�����Ս�t�+i��ݚ��#���Eֻ�j�ɦZdj�eTk�����=��+��.�ɧ,
b;�z���m�P�����K}�f�uD�=�s/ZW�T���P�{|rz��d���@6p��aե�B<�P@�P{w��������-1���2����SI���HGu�6�	���[y�HH�$;��E�T��P�q
�A�~bB�j���#�^��P	�V��*��>dJ.rx���:I%|	�|��׃�E}�]��wW�ލS���X߽)��a/cs ޏ��GH�j̹�|b�C��K��(B%�k�n�S#���z$�2!y�FBEC�JK�{@`�Xh��	 =rm3�GLe��DW讅�Yj���x#����l�6���	镛�f�v���YG�4$%�;��w������%�1G�nx���Q���h��8��d�bl?�Y<�r�0��
T���R�]Եm���j�R_�Q�m�3,>~vOQ��z4n4l;�obu����Ms��S���p0UZ��U7#����M������bՀh�?������}�'46�
�K+_kcj3og�]��������K��R�^��.������m���I�؛�,e��.���<W��Z2$������A/r;�Aj
��"�@{e:.��ob�M�S׀H���8��.�*�/���O0�'JQe�����G`��W�&�����R}��o9R�����4+a��O�%q�����P�%�g���n.��:qfȱ��`:z0�B�g��^��̚��Z6Z���\ �\(�z:��f������[��S�E��l�O�w���4R7�Z��g7�m=xa�7��8���U���wK?a��ql�_�� v���Z w.��橓C�C��ac�;���o𧻓׃�|H�3?�>�G�{ �X10�^L��C��Cɂ_���Ֆh9uɴ��C��<(����hm����Ѣo��p�E ���Z����)�G"�wZfǋ���p4kx_���D�3[�v��x�gh��d�9:a��8�oi�u���:��r��9S%X�8ťE����; Bz�<����G���zA㇕Ū)��hHe2�f�'���p
t$����|��w�n4?4�!=�ad��'U�-��dP�o#�l�XR{�}�"l�0c��>���a�����*���.!92*���y�*���%����q��z�̬�����@Fn����Z�ؤH���B�rDoԣ[U[�Hζ�6˸B�k�ɰ��,^�!{K䂏0�������E�������J�4>� aǷ��F-����w�o�	����~0Z�J�z}���V�fv��RUC����=9pE�)J��c�,7��Y���p�3SB���D�x�о��yi)�x����i���" ����\J�ڒ�Ѕl�{�c�U��VHޯ��	˽t?Vn+����jpzD�������x�S=�k���j���׮/2	���oQ=K!�lz/Ys}p} ��yp(����9?�MD�EF9���������q�L�HP��IK��G���r� ����q^v��8KP�DiJ;;����I]ߘs3������ ����mX�`1���|-o�Յu�7y��Xؤ�		7Uͤ��\��5.'�6���)��]��x"�U�be�S��W*��AI(���L�mq2/0!Nf����w�1�UR�9;S���~��	3[�}�(D��}�Q�����>�ו���
Y/\/L�o�p��n���p)i����*����� >w�A� l�,A�>9��\o0�� 1s�e�;!���*�D�m_;���	�ls���ϗ�@���U�ۛ9�b-�ܯ�<�i�%ԤRBaa�'Jd�g20�
i�Z��A3���������VOx�z[hjˢ��CA��bH��b�@�;2�����T�o��x��-p,lҾ	��n��a�U+c�@�~��f��hװ�R�z�}�>�ͅf2�rU�F�]X��[ܽ�[�C7�����p��������dV�K�����)0o�c3Z�Q/�Dz�;�8^M��U��Ӛ,��S�g*G"�g���2����P$ ���xWCʕ13�H��Gwu�n�������3�����\�]��ʗ]��r&K���5u̢`l�����m���ʹ��C����1+��FP��QR%�?WB��*�4;�>�=cGL��O�:���z�Z�(��Y�1����*��Ԇs5���\9T�5�;H���Guɕ+�����%ϖ8gH&1R��Q�2���?�ij«�Ǌ<V��,��q[�L$bj�����$WvO���� FK��
�?��53\-UaH�}�����C����F���(-s4���#�d��e�
:�V�"��\�9����h��P=��K������A���2�6l��F-�h�u����WZ�ka�5hR�對_F�W�i��:o���5X-�*_�P��?�
@�I�_#��IjZ��{J;˔;�bJ�Ko��������t'9j�� �e�xa&�=��'���kDZJ�?s�ª��&f�盱�d � �y�d�����b\P�W�',iӻ�hc�вף��(� R�G�0J��$��ٯ�2�^ڲ�=<SVa�8r�C�=�6c��a���ܚ.[(��8�����@�E����]���g�J`�ʞ�K^_6l�~� jx']K*5���]�z�}\`*,6�`������Ͻ�<ё[���x�͵H����,���\qP��SN�|���j!��&D߹��_}�?29�� %S-~M6�t��ȁ'tm{'0�f��:��	*�;(���\�j֟�Tؚ�Į�o��z�ӓLK� �yA��;)���6�C��?_G�
��u�g��w�����|m�~F��, �{:��N��|�ڟ�b���?i�ȫ9v4-����J�רLO|U�wN�B�S)�3n�'�~�潗>}o'��̲W+c��������b+y�3k��P0�p�pJ�՗���EZL�I��
���[>�@8���Cs��fA�˓�$ɺ��7q�'{���'�Yj�rq�sn�F��G�	��h!�$<�%����8Q�=�<���w�G�|t�� ���CjĐQf�	;Q���aZ:|��sr���Ǚ{��,肀鯛�o�T]����?�l��C������rV�q&92���8u��]�.��j�Q�d /n�Wk��m7�4"�X+�ũ<�y(o��9����=�&��"��yP��F�5B�x���9�1���Dkk��$��o����Ŀ�\�Zt�ƇQ:ԼyI�X�`i��]��%��"�.� |N��l>��^Na��!jH���I;�@�	)���4�՛d�	�L��x��9��R�ڜ\ޡ���t�<�~q��~�Pu����g������<���Y�Gz�I�\��Ԇgw�i\`aj;���<��Z�-�m��<��5J8,��}
�����!�0|S\ca�Iմ���V��M �P�KCu�=ّ4v �4rQ52���OraGd�-�j��)z�2���x���*C���h�]����	��+��I�^m]U�C��V�6�ZEVOpg�83!N�����R]5M@s9�����q�[ί�?ޠ:���4K��ᐥC|�d�ig�������zՊY�ߵ�m1y�/B�G�6�SL�n�i=�����PA�8�"1�30A��x�o�!�"-/�<S�ύ5��"�W�o�}�.#\u�F!��Lh-GC|�Cܟ���ݎ��2[��o(� ���7k�?fJp���V��a��C[����)h�
'�8�(؞�=L'�:�G6kh�-1�Ev�h��_�s�V��Q��&Q$���O"�h�;%����(.i�X��jf?ID�[���&.N���IeHwӃ;�M�:� ��<�"���]P��V��C]�*S��8xwh���zu=�3z�CR2�iW~� �L*���}�s�H&<�o���*�ǎ�lp)��-~Y걝��?�!�f�0ZK�߫P�D��z1��.�/ �2���q��2��I�$�h��-F�V_��J�f�'ܦ����{IC}���&������D�.��I���\A�P&�u��KPho��G9���C5	 4g%�!|�V����dB���˜
Vqy���d�f`!Ro�s�$�s
<z��?t�LN�w�w�W�[`�8�����Y�}�F����o�Xh #:�����5Q�NP1W���_�j�궨W8!�k��鸩�\Eo���j<�~9�&I�H�:6����y���UH�;͂
�Cշ�M[d�!I3E%��8�>�����8=o2+�y
@�(�jJ?�}�H{�4�Ap��/Q_A�v�V�.�	d��%Q]� �.d��G�K���#�K�='�<�UUՄs��D��!|\%��P�����E���J���)�HV����cE��"�>�#ED��"�y�ܐ
��r���5���Gq*�4�*�x��k��~��"kb0��Ԕ�}�["d���G8�3A3�+��9_("8X���������zo=��a��L�s���t�Z�D:���<���|�(���(Ֆ�[����+|D)c��.e)������!�-SxkE����n��g�����̥���*�;��G+�B�=�OZ}��)��/-��}�!���;�]�vîu�䜜��G
��N��tti[��PF��շ>e0>�^��'��z����aEC�2��RA�-W��`%!�_{��E��j?~
���W'�N���۟9�oKX��.�=F��C2����� w�%O�784|�޻0�ɪ]��	S��
g�Xw6��z�\/��)��~k?��-��84'{5h�@{2d���gEs��,����wT�����q�W��4wr�*]��ڹ��Yo.��ʏo���e��I��j/jK-1�Edȫ�e�rK��B�X�6����@� �kκ~�\	���a0ȋ�hm��=X�+؅���X� 7[EjC!� ��5���؟�.������ |3$B�o�&���r�)����L1i|3��g߁���#�-�H�1�|�K'��LG˴D���&�=�t���\�ԩ.Z��ew�0��Z�������E#k�RPZ+�&Ty4{u��Pn�:��{_ ���+������Hm��d.bTfV0� ����<?�4ږP�����4u�ra����f7���ڰ�^��3���:x"d�3äOU����c3j�@���0�ma�� ��Q4s�V���%�P���F����N��PI*����a]/٧Ob���VD(�}���k����b��:\,��ߙQ?6/g�	����P�5�&�2�h��ng���={�r+m�lD;�F�{xB@�W9��BD����*�C�*u�Bu�܇NL��6��637J�`u��p��R 4,�*X)/Y/�ity ����t%#���k�D�Е���k�'���?{��F��E��rn��)v6�l�B�\<2��&�;��gk�<]����E�P��zѵr�8f�������������&��JO�N�(�{&�������P1j����V�%E+�uU�zM�^_0B�).<�I)���ğ��8�뵹�N\3�!>o����N�a�S`�᥉Eۨ��f�\�4��8��]����/<�����uh�Y"��Jm<�Ps��"1��@qp���͛ح�������/����!<��ry$�fv�1*�����_6x>��N�%��+�z�� ��?�:�6�PLa5.��W�x�z�[V0�"zD�Ȇ�c,ɐH̖��A����?���ج�ʱ>6?�U����{��-d{�g��j�Y�K��W��%I�5��`���Nen�J*�FJ�t@a�����,��^����ݢҟ6��4�;b��WTQ�i<;����W|�T�"u_�i8,7u��[tF6��H�e�YA��1.}J��j����{�LH �eB�6�"���B"'��M�aaY`�྄. ��%#keO_s���"����\�<:�3'��@P�ݡ{v�վY�J �᧬�L�U���������N~i�CP�:hYH� E�a��7���=yH�o(˾E��{-�Dl9>�
[e����<��V�Y3�Z�47�{����yT@m��i!V<�m6j�`�=�KL7hB�S�1?%��hW%5m�K��4�����IA��ۦ��5�"R�j��9�2��<ɑY������_��<���E�l���3q�+CuZ����I�@� N�%�����}^88�S���Y�� P�q��q�0�=�d��JTB����:��Wn�Cm�w����*k��+�F�
�"�@b}]���SzJ�������RN-��D�Nl���V���b���D�q��j.�W1׿�}��`�:�F������S�1���ZO��:���u�����A|�!������xQI�S.�0�O�I�ٲ7.V[��a��bmk�Z�����-V�T"�^�Z�ѫ�E�r�ku�P�nA�p|\i�2{m������툮���0s,���iЋ�YhB�;()���	am3�U�ص3ӁAOt�,� ��bG�4���E�������5���Y:�&�5�D����!��5����=z�o�������=��Q(_��O���ISC?|�z�nɉ�$<�~�f$�L�u/pZbYs@U�|S~���f�
��
��H����}�?�rW�|G G:�m�tD�#��w*=7�{�O1�#���"�����ƌ_���T�=��B�r6��o�6~㛴����!h�i��֌T�_������b����(G��"����/`B��w��1�H9�^Z�I��D����`�o���.�$��
jψ{/��uR�9��'GQ.& �*�q������˟�@9M��O����s�ϴ֏.3Y^p�!S��+��R�j��5*� �E���2M�J�����235u>�CE����f�G��oK����CPfh����Ѳ����P����'s���Ӽ�K�ؠƊ
CG�@���.�����v�8q���\��s*��|3R��0�4�6����
��Ğ�P,6�%�3_�#��Q#���|Y��؂;戕�$s;'��)�	��蟤���]%Wz�0"@�P��Gds�GFQ���������T��/�b\����J�0�v̊�0��H��:@K����y��E!�Qt��t*
ihMk�Ø���`+/��!,��^���� t�5�ʠ�=�ЇH"�����(�X+���4�0/5�F����-u��<����%Vy��KЛ��+��re#U��:��7On��x�����?z;qXS-�~:^��(��[���[�LMΨ-���;&�0{6����-e���Qu�g�J����w&�K-Ț�D�/�S�׬��'���?�)jX���Q��)MK��f��!x���P�]�8Ft+�1��H�(��
5�� �Ri��N�r4FB����R����nS��jy~�.y��\���i�	v�>y���8�~����\�u��z]I[U�����e�va�fP�ů[�<%%����M_ـ���$Ek�4Z2Ί�����;��j�l_t�<�B�m�c�1>�LQ��TEA-��LP����rF�T v˒�� (
�B��r�L�w�.���=Y��~�6*����%�[tFKfp+Æ)�<���\��	����(�b���b�� ��g�Meg�+��=I�G��qJ<G����;{�0�����
��1��`��ꯂW1���>����(~�i1 �k`�pO]����FaM����3����He���_����.$����
����v��e��ڰ�;w{�4����1��D��f(Rv�I�P��;�C:�㞻��K��/9(g	�(L�e�(}6}�Ѷ£:�>i��X:ԋ	M����C1䯄Obd6�c�.8��a;�D��z���)5����W[x�-�Rʎ��C@����^����ej��Z�٢rI��-�����jcr�W�ꕇ�Wܙ���������L�ػ�w÷��&�CNl:�JV=��	��
�(i/���]X�X�NKqGS����pd�s��[�-�Sf۲c�,���f�U֦��_��[�EfOt�j,��j�Sƭ�K�e9�u�B�[�m��2��t߶��xw� p	�MҚ�;n�n����z�㽌=w�E7��ڵ{�I������!�"��v?;�2�ER��l����	T pjȭ�~�K�*����z�n/P�¾�eq�##��j3@�ܭ|M���Ҁ8G/γ,R����YZ������"�ۏ�4i�6Lzʰ�(��������nA\������p��ץGaK�B�h�D��D�WF��{̝����zj6 [���)U��Z��P��'�9:�";����!{mr��/�iP��\�����N���`���P-�G3���`~���L�tN�E��f,P���ą�9�$k� �6�l|k���vr�1���v�?y���X�����ڹ[��[r�S<�F(2�݊jþݠ�����!�Ł3��x�㦿���x�R����f�Ov;�9���L�R��A>T5r��傮�9�gʶ�'��&L�0�����|'����m=�gw]��h���h�H�ĆؒH���<\1,
t$n�`$r���(҃���nA���vE��Z��j�����CX� �F���Um"�ͨ�H"��M&8٭�)n�k8����~�Ԑ�x
�w�~���� ͷ���J���%�V�/���B�iYf�wL�~#��@�S���NXa����4����U��f(?֫򘨝i�&9�td����ץ7t�.?fm-MܲHj~jXG-��,��/�$}l7�z׍��hD;&�3�ey](2�(���g�ܟ�u/Oљ��9%�n�g��l�k���	�����q/�)��0� � a<�(D�Ma��Oo�5A7����ئ>���� �����'���qo���M*s��� Í�Q
s��i�&��eӺ��h�p�dn�wLt��G�D�6l~r�0�����p*h���"���(_{
o��Cc%����'���Ae��r�zE"�cΰR3�Z<Һ}����_\�{��KŞ��ũ����o���;������`p
���dD�9�o
dS/�Q�@~�O[�ꨊ��6�[#�?|I<���S�G^�_\�8������5U4L�!�T1a89;��	����F�LhD�8
+
�[���q[{�h�fsxܠ��;HA��e�1������#z3��}��ߘ�ǿ��_Y���a2����Tɝ��[E4%��Ow��W6�ɫuh# �u��,��
�`����!dd�.&�j99?i\��v搜�kЋ�`{J2��kD����4��w�A�~0hD��H�ć���u|Z<TzP���	������Qh��q!G��鏉�0T�1�\��;F4 �����QzXwz�l�h�q�:H�@U��h�!rRGo���E�ɭ���?�`�y)H4L���c����ʞ���_l�O*������-�S5�93/��bsE�ӻsSLM�j�:@�_�<r���. [��Gh��R��5]�O�B�����`_ӏ{�d[NE�[X������-?��`�*���	�4����w��SYh;\�����hۇ���c�'Nupe� 9e�ke<mUQ�����8�Zv"AȬ�c���_���5��3�8�QN�J��M(�a3ߘ�}DAMH0�o�����A�ӛ��f ,��9��g6nyK��_�M$��[�s���qPqa���Z����z����(�&ŕ�/�Y�?cĤkR��R�f�q� 8_�f���"��Ȣ���/O���[[�oT��$�M�(�>f����z �ǆmO2Z���h�[�#y�g���en�4�K3x�[�דB]��ɧ���h��z;���(�	�������`����=��A4{,����]�'�����ٙ�t��*B���4�WZ̛h:�k ���� V��s�w��2��U�xK$(���4��zVI���R��v�ȑ� �8�\��B�j\����b߮�'�����u
	,<ǋ���	��p<%���z�[?;�!�!��^G��c���Lt�8J>�,�d����r��VN�~} ���E�p�i� �g��O���u-zu0/�����v>��<r�����9�P��)�����*���t�@-j<�/2�[�×�1�(H��XJ�&a$)��$�D0G@d�t����-�t��k�"���;LU�/����FB�2�n�HJ:EB�#KϾ9���<1~RJx8�;�椄
�%��	v.�2����^�%N�'Y�u���q5��\Ne�b�G"���_�>�RR��5�{P�N�I�w�Gb,�E��g%��ؼ����7�'�G��FΡ�}�R8�YW5<a�E/ؼ�>����x>�?�"	��~��$����z*}��4�AEf�%� �H��-���]m�^�m�:��O-"ujj:�i�k��:��X9��b��1Wc�vd�����h��Y%�6��5��Xb�8�Ů)��C�N��A�Z��?�*�L�"��s�Q�K 6��~&.�>��
{ L�����ߨ�9���Q�	��������I��k�\l]�)xP�g����?��W����&����������+z��#�n[���jZ۲n1稏ӭޜZ�'P�R�vD���ro�����:���S� U��!gLd�;��v�$�G�p��[\`���_WQ�Y%jJ�f ^m�_HH�p&p��g��j#����K��
!�V`d\u� �I�=�UG�ˎ���uq�1CPsO��.��ٱ�	���?��O����r?��u�޴l�k�O5��z���A&�CX�Q@�����H6���qՓ6r+��_	n#i��9K[	4�;�^[�����Æ���wzR2x��q���.����Q��o�dwZ4���v4�柷A�/�6k���ww�@�hԅo������e�l��a�(�A�	�6����;�u��C������y�)�ޓPM��͝�Qƕ�`Sϣ�*�U"!�>���c��P�;�{�_Ā/L�^j�G���fƐ��t!����/�3���'h����yqaį��9��<C'��n��W�1�� �i�"�P�<��zd�X�d2F����JAM5v�6:v}Q�Q�e[��T���h݅�1_Yj2:� Ϧ������5�*�$�S�o�Kӏ��Ix�(�*5��a;GBUz��n�A�����n��i�L�����v�♹"k-�'5Tp6�鮫���� ��=rg�4���s�I_���Jʪj��'�{r��j��Yt�+O�Wl���_U��-<�Nc���%��kQ�w�!x*w�oP�QmU"N-�cq`5�_�%���S�)@����Ҋ5���[h�x;[�;�j)��������r"s�<�`<��E�6-sޟ,8�RqK�e��%��
W���:��	<�~�{��.�m��S~`�x��N���D�tr�=B���T7�ʔ'[ퟻ���M�@K+���z�v)�Óp�]Ŵ���|��!p��l�[Ie3׌Fw�ك\���3!V���9[� x�d�b�P����������(�R~対����=a�9m�[�o:Q4�qa�6���D�ȤZ�L��:)�׍�ͺ�S͝*�w�I��0a.����l�^�vy�	���OI��í�\h���>�V����3*�Q���<�_S$�ȓxS��Y1`ow�<��҇xJ�uć$�S�s���XK1VϛQ�r ��T5��d����9w�X�Ɣh^,�_��'}���9s�(<e	��~e�����U�Av[<~8���s�����~�vgQ����������a���(vy�������"���~RR8���J��{�)��k�s���E?�l���̂ô�'D�� #`��H��1�}BbJ�u:�P)��@�:j{�ݪ���aq�F�#�t����#�sY��2¡lxEVK.�I���U+?:� �?����T�0ń
����~�Y�87�*���R���mB���S�t-���c���*��p@ o}�9T�	�@�:�fZ�v��%^X�[�5���������5�;G5f��Ɔ���F��� ~�J1��sz��!���~���k[<��%̧�|#+���"f�p_�![b�D�}�`Z�����4Dn�t*�r�f�7�=j	W���U��#m����5��A���:��\�UC`����8-���![T�b�P�&n; +�n���U� �ܽ���;s��2���-�O�Z��CSF��A���IEۉ[�1W��<�8^h�5��^�3��2�L�����3R�65���Kć���:�9܌�BᆅEp�8V�Os1�c��2ݮ�ECԦqN�USP��<-ۆ`w�l�a	���������H \�Q��N~4`DX��s�`	�2W�N�6*9򉤅`�Ἳ)Rl���Ģ^�&��˕�|zd?	��V�#����Pc7�6Ń��R�G�h�|ʀ�x	�Y��D�8�Gv���lBf��^���{��9����r�4Z�Ϡ�?30�?$�J�+�t��G�ړ�h��#��>����<�� �W+��ſM�0��b�{����AH����Q��W��|���]�%�UE{49�L[�zד�pA<�S�.Q��TqCA�]WjT�+J�� }j�iS�!x�B^�>�psv�0#Dzf�0�w���w[�pNq~(���q����Q0VR���qy&Rd�in8_�G���(�쯪�ʹp� �(���q:x+EM����՚�Hf&����+cL5�Jv��zL0��z�%���Y��e���{��S�������B7m� �,St���G/��G{�(�0��$�b�1���ח��:O�������<'cY�F���cq���Y����:_�$��������LW���Q�fq��Q�7�����c�EF�i	��^�jy�M/y-�DlT��n���F�3���S5�*?��6/�c�a��AK&���G��"_�B��Y��1N�T�nS9^g�����9%�����~2+)߲#oFYs�`$�M�!*�K��S������6��r�=�,��U��~�0���gb�R�P� ����WIc�D>�s"~4z��$��� 7�_���W��'zVO���]۷K��ԯ2��lr{���6B��l���߮����|�k��*;�8�x�.{�A�ʢ=��@�|'�"�c�)��	p5�b&�1	;�P9&
����o�pa�qf��k0;��0���:�K�Y�#�X�&�s4[v���_\	��=�0���0͍{��l�TF���P��݃yD8pk毡`��� ٴ]C�
�b�6�A�l+�u+�!�|VIk�>��J /4T�2(���1���vԈZq�� �rQ*�kl��T�K�Ǵ�]�S��y��t:Zr>�� �_4c����w�0E�ߏ��?O���U��n0Ƙo��w����J�QO��Y��
�H�ӗϱ�șf)��\+����qiQ�o�گ� fʔ�4��۫��㤜#�{� `���cSͼ#���iu�"-\8_d���^R(X[�D����FH�'>��C3�<�f׫t�÷uM�ǩ�)���2�)}h�����@�����$Eq����H#^�T�0��p����ܸ�"�׼��Ì�q�V߈. X���،$٣��1]D��kn�%4�:�(���������;���P�:?:���{�V���L����'m���Z��7�B,��
�kN��a��΋���[]�H@�D�aD%8�%���w@t*��.�Ͽ��'�/�Z�'�W=A�������\+�ìD��3��H�@G�Eh4G=����r�N��V�}��y5��:%Y{<a��M�*��/�D?U��V����ơVff�у�B��A�)���`zdQdҁ��e�e;)'ۉn�/��"� @�B{ƅ1vmF'�͛�(��B4��{�<�����bj~gўn%��[4�%��m�v>v�q�w4lL!�f�w�^
w���wK�]
%�V��R��Y׶��Gϟ-�vY�Y6+�[P��=K��ךH�������������W�iܿ|�9���y�H��{$��
��n��4�F�g�(|`����I[��4�#;�U ����O0��a^���%�I`��+�dZ��4PnB�c�ɩ����Nl�����o)���k���p���}����h#e���1{� mH��'���,6<���`ok�W�9c����Ɇ��Xmw�NEl6%�\R�=�f�<����.ફ�u����S꧄UX3��Ķ��n��~�	��T�����%��	FU�����;�Q��ܷ�+�4��QUӲQm���:��?;O�X},�p_�f��X�W�̑�m�4�'ž���_�����5��G���PQ����v�����i���+��K%���g��z�
�H9��/��n:��dK.2J`s��LGQ����wK�[y�qނ��>�q�	��%�G�iS�<��$�44��dX�K����V����J_9-{�Мg���g� �_^Y�.�f�ʏ�_$Y��Y�1�f���^�xJ�^33�(����f�7�*��De�d�4�JK���+.�e�T����A������j�_*�d�2�fz��V:~�po�rn�N��{$K�����i��3ɋښ�j�V�b�q��g�j
�|�v�FLb�l�>��_��]�V�F��):�0�fi����i���e��n�m�
��h|�����NkR��W�+�^��hK�ep�P�B�M������>�26.3�#�^4��V��a�k�������H��7�v[d���P	<���W%���]ү�)k,���|��g���H�P(����H��{Y-�+��4 Z�����.����%���2��N0�#{��ް���^/(�{���ȝr%rǑK�e� ���B���/��S�t�Q��Z ��tk}��-x1���-�?"\��Wf�^4n蒫��m'�^
E٣R��F�&���%��K?��J|���]:-�4�K��tH|VuR�?]��g�c�=a����uU���)kNϩ�V�n�{��:9s/d�pV�1��V�A^���Ί&g0tv�P�-���l��'����.ߵu��0}Z��)@]��jYN�2RR��*��dxPo5�4����S�ٕ���|�UH��0X����3���C�q�$&�Gq᧍JQ>/yfcJ� g���Of)/ϗX*�*fWt���#?%Ͽ?oRc�I��� ^(�c��Vrm>҈_��z�6��!���B�����y9����^��,��<�-_�l���n���$<>ךD�$�4W��������8�h�6��Z;g�VY,������d�w�5�&z͏a߼Gh�z�*�H�$@�8'��5��$޵4i�l�W-��J�ׇ�$�YG:/������;���&!�0
�꺴�[�U�1�ކ��zb�ݮ��e�6�{�i�_�0��Q���k(C�K���D�I	���ͭ1�/����I��U�&����${�I�S���rξS+L&~���#��������}k�z`���I#�,��&��ܹ!V�5�ihq/�D���F�?�B �<��(��M�pb��ah�)�ё�dc�v(�1�s�f��C������"./z̦'���k�(ǜ�1�n��(�2x�cG9���i5��J�����Y,�2s�PU�䮡���U��9e=m@[��
�`Rkg��� j�dڞ9Tm62��3�TL��W^{�2J��2V����5 JѾ���Z ��qanH����9+&����z.#��l��To$r*,�[��vq����r��1�2� ���Ш�(�\�{ӥ�"7U��C�p�toi��̟/�to	r�1�un����V(�v��4�@�)�?�mSv�DTQۓ%�.���6�n��Wr�p�����t��W���#���S���8NV��=qf���zc��s���F��p���u�uF>�ؠB=WB�&&���(e���� U�f��'� V~m	�X?\�{�M��zP�#�VW�m:Gd~�i_,�׾u^A7�����,�/���'q�he&���U��,�.*#�N$n�#�-����?��MQ1��Kf�%*a�=�i�T���m�}L9Ӏ{�V�G%���B(r��L����;�Y��-��&�>�甶P�ҖFg�?��n��zW�3^=�K(� ,�+�]�R�V��X+�K�I�i����Cr�a��eω���fQ�Ҍ��N�<��M�"LE��j��	8�):�_1{P�^�"����&�7S�@�+6�s/�+�G�W�l�_r�\"�CΤ7�Ѣ7�T��A`��#&6��;&�f._ y.�h^>,�)�+t@;S�_�F��i@@�]�JD�'xs��۽o��M�&*��B$$:4��H?]��o.���n��BP�Vn�斖�^���sݒ�r��˘��Hq4���z�d�#p~Ӫ��>P��F��6����x��3�}{ Kj�%p+�h}��+�6A�����%�H��%�����"#O|}�O��g���v�}~a܅��ٞ[�'5r�@��y⾮�1	��!}8���߷n�s��6q����ƚ���m���b�j�}��U���D�q��� ��� حuR�6J�-���8�a�\��Y�K+f���D�{��u ����2j�E�r�ou�WN^����,���;H���ƕ�ʬ��	�a���D��� ��2��L�*X��[b�(I��;F޾��T����-); �`���#z�8F�q��+?H�IBU��#qY0����!�t�D^o6*E&5 Y#�j/0�gh�a�)�&��+�#�0z}^v<�xܹq`��]W�DP2�SlM�2�+���b�G<|�k��:�-bam�W��dQ���Ɯ���N"(|��((�j�"�)e�U�g\��o�Jh�73ϒ!�iAk��+%l�N\\��H�l��+���Ue�h��z[��ֶ����T��z�d!6����M�p7S=�p4��-��ɹ�ˇ�f�~��W��6��"��Y�B����W��x��Qr	v6D����-�G��/`�	y?ؾ�� X���(��D��N��Z��Er cZ���DX����`����t
X��`1�I��6P;�c�M5��o|������r�%ܚ�QЭ�?Z�h�{��Y�?y��Z���iU��^g����r� E�=���g[��_^�� �b��~Sq�#�P�u��O��xIdZU��E�!�O� ʧzK�P�2��|3_z���;Tza�y��{_eb���߉�ht�Ek�#�d���&@	g�aԋPG�ļ.���*=��b��'66��T^I������LmB��Q�Y5��xgН@�Y30�y�#�^���N�[x���,��c@1��+�+ʕ�K�GVs(�����0�����a�@����L�~9�����UL -�ϫ�]�-��s�\������maU�dE��JՀJ*�c86�R���oq��3�C$���W2� B�����V��v��c��D�}����ٔN���@��K����p�]_�7�����E�)��W�U�i7XE-\򳋖4]$�=J��Y���&Ӽ��\��oe9aSgH����t֋�������l/{C���$���y��*��HR�~H���6�w�(�N��3�l/��z�#��8��V��*��q䛸��k��r��Uy4)�:��d��"dK�zǔ�ͳ��r����OB��LPy�WHQ�j�RBA��B��jl�tÚ(��A��W����/�W\k�z��%�%�� zi��b��C�"Cp�F�����2��<� v� �cG<�	�V�Ed/H�&H4^���rF�%-*/�!+��A�u)Sg��S�$���#䔀�k�pU�0pp������w�����1��n���
#sޯkq~�FU���}��Z@S��"�^uzEf�l���x����X���YmZ4�o��ݟf���a�-oU��W��Oh��y>�Cn�ߒ�5�W�S�T�}2���kI�N	�={�L�`��3*�0����h^�zZ�QXa�y����	O�*T�l�8�XL
�$��v��*��$ٺXD���i�s��ɡ6z_�s�2P��qCjK��f���	�7J����3�[��U�,%y�V�/f�y�
1�!�>ѷ�E���_5��cj2�?	r���P�$߸��� �r����)�]���s��Ϝs=���s��W�F�#�R�B�����V�&�w�1�u���F�K���Bo��S^����VN �}n<
�v ��5�����R����H
i�G��s�ݢ�GUp�� b�$���?۔�;-Hu@����O 8��m&�oӷ��t8��&���+�?�H:y#��EN��p�1�r�;q;Yh?Piʗ��`�KV+$^��V����K�[���*֟�5R��Eӓ)�qP[�1���b?���P�
r����?�����(�T&�����y�(r���{T�_jF(��iY*���sXf)�⚖7
����:Մ)^Y���-^�B�����= �T�`*�y; C�цX���K@�8F���#G���;YT6�S�,��4y����_�ƁM8z����z�S @��a��ݙ�[I �L��/��R�s���d�"؜�7����^h[�y�;t�-�x�2�ځ�c�����@�G�k�dq=�W��T��� �C�#9�J��]č��n��9R/���u.n��[�:�p��D�:�[����%���|w�U���2�"�"zu�G٩A2���7���q?N���O�9q�`�%���M�V-�`�B��OmӉ�i]�����LLfѐG�n�M���n�j����s.݅���� {�0qB͚��mI�_&Gٜ����o�6�n�T���1��wW�s��"w0��-}
�_��h5I�*E��� }4ҝ}���|jr#+a��/hA��6�
�{ŨX�Ӡ�I�������tL,Gz���V�uو�D˧�7E�?�Xa���@�Sw�V⺬��]r:�D?e�]��n߬퉒%����:&��/{=��h����*S��"�*�ih��h�ݪ0�g3si2�k�/1����DE!J��l��j�p$t*�M��wrg�����%]��t3��?��B� ����8
�̂J�eo/�z��[1�dC$#Q��PRI��'�p  M��\F�m�rL���Z'82y<|	wp��țJ-۾J7��:���&R�y6��z1C�#JP�q󞯆��y���`�&���)��7���l�[qt���-��<%�J��E�/K^ĝ�_AB���g���`��oN�UL�|�~�;W�v{u��	n���N�ڞ���熆�Vi��	,)8S1�Hwq���Z~�����T��1�!��k��>�?�%��{�Ú�@;myw8�����r���-����[i�V���X�
=��K�����h�VjodY�j����j���uW��Y��Y�0�� ��"���p�D�4Q�`�@�r��sI�^'J�{��+A��h��,������J�5`�k��	�[���PBX�c�Ƅ��x|����J���|\� ��^)���eنS�HW!k�M�j�8/��6V[�X�%���Ο�-�{C~y?h��Ԫ����B�i�(B���ɚj���䦧��,!Ack����F==L���L�7��gg9�yN��)�gE���}N�
�9��	��5d��X���H��|���^�嫩��
���']ng)�X��7O��|KĻ���5��~� �UeY�����O�DԐVQ��Դ���ңJC�G��� �)��bC��P�G(zV��$c^`��>���I]�-��u����o?���@wӐ�Un�r5xlC,�"�
��Qc��l��K�Pw0��y�y73��p?Op2M�����,� ��L,�Z���uV���a@�֎ԡ�qnN:�#��0j�"�j��R�yeidg̮��SU�ʔ�d�J�o��1�в�$�GU���[.�tg��W��c��e|���`��&~�O)��6.�+�V�FjC��:I'��
y8����.�JћO�H��'+�2��_��R�A0!)�7��0NGԹ�P�iG�QH�TD���?�L�i�n�k�z��8Ȫ��oP7x���5�w�kw9��7�LiݧѢ9O��%.Jހ�|����=��C�M��T��w�����͐�����c��U�P=G3#~.0�8ܝW_��H�풐�'�5o8lъM�[G:�L������/h,�~]��l���L�{B�߲�^�ȳF5	�C�M���Jۭ�"���߼t+I�~�[�0�${m�kҸ=�R�B-ɱ���ڤD*�������j6�k�Ũv�ʸ�8ÔnuX����SP��ׯ=��xM�c���l�5���l����.�G�4���)��p� �����g���� �'�G�Bz�WK���Bh����� y��YІ��c�R�줎�Fh$#ހ�*���;���K�!]6�\�rG?�Zf��Z-���S������-�&I�Ù��8M�{C8XzY������QU&�E�D�U36�ٿ>�8���/�����	}��8�
���ئ���a��[��Y�ܲ_���U�B?z�YoW�)#�݀^)�w�1�='z�+gӀ�!K!(oi��*WDRSq�E���$��4����8����У7��M�;k���ʾ ���y9L{�.��2�8�=���_a���'�-毇��&�ǡ>��
�	��Z3�T�]�x�v�+�
�-QA�A�t�r�B��������&�j��r���G��Hj�.���p�{ӷx�-�_�!�=�tm�W@�|!n8�&��0L�J�KH\}���N��N�Jz���~�Rʢp x0�W�$?�v*�%��Η��ͺ*�4�������]Bv��-,�������H�$����^�gq+U��r8m� �(���C�?�^�3[��n��;R��S�����/e��L����V����p��T�swh�����L�,����k�a�<��"d�p���tOԝ��1v��_
H}��I�1V_�ײ����M�U긑��y�z�ֈ}d,^����u����@�+���q��e�	̲�-�}�U�(��֩�6�4'�&�^;�s�ϓ�Ŋ�:5vɢu��p<a~[;����4p�gټ����/c�B*}�Ó�OkB��Ʊ�L)ǂ�^��E�ϙF�x�(��e��)���f
U΅�ld��sԤof�?�8d�@� ��V��J��Pl��߄SO-�9?G9�tJ\�IX;W65U�uU'�o�B��W�W2[s��o��'����b��yB���r�N^7���eߞ��fM�uVy�Y�N;�/��|@%�QJ�,'B��e[$�p����]H�n�x�Ǒ��?�J�d��R�*7 ��N�gòT���0B��m{��b~�K�x˭"�Q7TR	Å�Y��4���ԗ$b�����%��&���	O�0�Z�! ?B=��	&��Ɲ�Ŏ`Ҵ`&�w���WC������)�i�D��!�-�t��V٢�bV?OE0Ұ9�ڊ[��N>?*11~gߝ�O8uI������1]��<=/�]q��XՇ��U�-�o��݀��b!"m�+�b�mWŸ�a9��.�:h�`;���C6�d-Ra��j���U������P"�gH���z\�L�P�'��1|0Wʠ����v��A�����b^��^(T-\y;k�ܱ1z1��om~�'W<�.��:��x��s���ő=C�C����	�#ae��|[Ho�I�Jt�+ʦ�;����z���S|��k��(�N����	��4&�B﹊r�]*A-�}�&@U�8�uS�T�1w:�B4�!O�x��rd��캏��d����1Z0�9g(Dx��� �Ʒ��������9��\���Cn���q��
2м`:cx�o��I��|�2:� �V���[�ַ�Q4���04>$�w��i�t�K��p�|�\�
�W���S���,��}}����j]��n'�D�Q'.<�Fr��?3=����efݏ��}���V 6 ���}�Rz$%��.h�(s/-��^�����TJ~��x[�d���5uK����(�K�H����#�'��ACk e˫���<O��l.�P1�@]���Xj�W�P�����G��R!�T��#��2��g��!g�m�U~���:-��->���΍'r��qn &9:#K�iT?���Gf���o8�u8*��)�h�4މ��k0Oi-�*�A��C�l��!V��#�U���6�t�R�r�5Q�๏Np��_a�/� ˸�Q2�aM�g��p^�U��ǒEtR�����_9��'��<LĈԲ��g��U�Q�����=�0)�T��BF1���#��!�t�uH|�63� 
0���>��_# B/1��r�wW<ç�ĵ=��_��Fq�@n�+�Աa)w��RF!����pح(*Aދ��m��n�װ��@�]�A!f�}��,|�A�Tu�� W���i����Ҏ4��R�X��(� ����O��)0����__O�NW�
cW6��h�^��7�n������G,�s��$�V�xE���/J�R�v�A�Z��4!ȧ�Y'����4�ua����왇�����7Vj�9�����^�(�5Lk	��~3�GGE���j	_��6���T�4s����/e����.���9i��7�����ւA��,�:��:��Tm܏���?z?�XU
�$5eKjGP!�2������]�@c�����GD���0�Eo�Zuc�xg>+qJ.�zތ}����5w(c�8�W��~Ę��D���h��!�5иy�u�m���,S-I���C0+ �ܿnq�fT8�]c~���o����<�sv&?�;Ԏ~�VR�V*$�����	��g�q�Ƽ��BuQ�*�
��o�V���L�t?��@���	Ki�e^�R0�X����Fwǵ�U���>�����ǵ��jrF�k�X�9��NN�C65@Sn��* (UF��x��V���O�g�n^J�� n<a����ŅRpfe�PR���B�M$�+���c���a?._�<V��Eqe�F�kA��;n���r���~�1�c�mH��2�O��O��F���|��_�=����ly�����"s�PI�
Ip�0KV^aO@Q���摬�pu���3Xji��ޥ_a��5Ѱ⾢U�u����+a�ev�*�ʱ���^���p�*�_l��F������´͟��!* �\Աe���E����^D�I�)���U1�q��W<��w�	z�F��;!�|���^�֥�0�Tl��l�����v�ZF��G�D�����_P�:�#�w�R,���)5�/ɶ�5l�*M�̖�b�^F-����dV2�SO���p`�<�3z���Ur�t4��.{h��1ᇤ�ܥs�2��&P� E����dT9��,�Tӆ0!��PO���.��s�=���-39����)��w/#�%v�ʫ�|`[�>Mշ�)7uʗ��G΋�ye�2�U�7�^�fc:N�E�q�jt2򰲊��$�7���8^��Q�3�F�hF�2o4H��0�e�=��ElU�,)I
�Ȗ`�Q������b�*;�~e�֙(��ծ77�;$? �q�c��(!&RL��t�j�n���a���+# B�=���a�H���@'9oSs2����
1`������Z�OS�����;��>���©�X�V�ʄ8�*���Y�6�i��
��1"WXÙ���#,��!�k����WCvR3�|�Az����CScLh�`u6=�B���z�d�؅9��R_��Jj'CbK�q�"zO?�i����;�L�o�:�{ �bX��`r�B�RM&�t^X���/_��)����:e�uZ��4�09I�=�?����@m��nN���N�-_�(���1.lv݌�{��i'M����K�rJ��ΛI�W��]"���	�8gχ}�i�n�
����$�CA�b�9&�/P��������ٞ�ё9!E�{�\)�7��|7"B���x0�-�Ǥ9||/ɏ�(ZFP���#g�l�?�tT- ����.�`���w�Mh%2!��Ou��0"�5�C6�n���e�P��o�.M������y�Jyz��!쎺�@#�"$��!v(��=��O�J����*������^)��BNF#��/,iR��/�Wٙ~�nypT|�+{��e~�����!v�I��Q(��v���_z���j�� �:�E�u�(D�[ȅf�?�!;X���{d�A2f��G~Y��c�i ����`�~]N=GzFf��a��dr�B�v.`S��ϰr��I ��_�TJm�ð�Koߜ��8��a���B2CH���2Q���D.�-'�P�����2'(�U�O|��>_������*l�W�*w6��{��G�[�<dR'���s`��0�֊gT�Sf9�7P���k�\����3�d!ҭӼ�#E4�ʾ�R�w/])�567W��A���@�a�5꘳�j�<��#�G�mU�=���!��L'ռ�-`xNc��k������!����_v?E�iY��O�:�,1v�����Gp��wc�\h�J<�Sg �w��1؊HJ:�>�A�1����e��P�Q��Q;��TC�[FV�e}�e���`�e��_��O?_���v&(L�&��#��C-��r��
t���vp l,��S��O ����g�YPa�X���>��F}�&���~�i����8�#*�VփRҷb_���\���{٧j~�]��8H[�DE�?0���Ֆ����y?����,��5�Cz��C�;J��ϓ��s�-Fv�j�{e�����ҭW�b!�^O�Z4KħQ��-ZY
hGq`U��h'HoVE fLhs�`��P2�^O,ݚt\,61j���S��g�&���y��Yv$	��r�\�X��1���0�dY� `�>�qY���~*���8�5��Ys���}~�[��Ei�����(�O2\i�}fQ��T��*��F1�:�p��$���M�?zd'�A\\݇�}$�,!I�^]M:ӭ�����)�j��@�J�d;�F17���N'��6��d��Q;K/�Ԧ`��u�']�_�s�#��/���G���*H4���b���(�^pуw�y��Ɂl�#m�X���hAm��)P�0B�P'V�O1�h;�{�U`I<���Z��k�bI]�ä��K���?O&/>	H�s���
:Pó���-�'K,�`�QA�K��Uo���/��q�"�(#���I�z�B�@�u�3�b\{�O���!��vF�},�.���?	�
����cK�jK�Q���/�b	Hn7�6>z���1Tմ$��)�3��� .~Ȝ�( ��g�?�8�Ϛ�0��_��u��j�
!E]��d���!1�b���J�.���8���vZ�pl�[�K�Z0�Sl��R�7�� αL��e(��~0\8�'��[��?����- {M��}K�|g��"��45c8�y�Q?�d�O~��S�[#q6�]�9�����,<&�O��"�Z�|�tz���O��#�#�H�0��6�a����Zk햏i��G(�u��~:�_��6�g��x�Q�S��w��q�r��R^�&+����ހLlPĈ���ί���}�o�Q ҷ�5'������M�ۏ& �I]4���5���z��NW #���O����[�r���I?��,ӗ�5��D5�ǇHr�*�u�"��4�j?h}rssyRgA��U�O�_y���p��.y�G\sݘ����C4�1��-�l��.5��iEZ�C�>�,�ro��g��$FÃf'��%v��@yb�@��rZr���c8iO��z3%���|��6�6��a�#�^:���P��(`���h�k�	_�JB��*�o���u���AW�@Xܜ���`�'l�|�����j~1�[�3G�N��JC��AVM%������ �nQ^Us���f�S%�Fԩ>t�PL�¼�!<V�*h�h0��؄�+�aRz�*e]�:���w�6.�>2L�Y�Ѓ�N�d��D�Z-�d�sG�Jg�Ƒ�BeT3��{�JCd>hf�+��0~j/�t�-�2> ��Lr���Ȭ�a6g����&,������+��1��gd.d��Wyp,r�th���Ԉ��4O�m
z�^�h�v�wwj;Ҥ�Z}������CQ���Q橈�͉Q٬�fPL!z�T�T���dW�	��2k3���Q6��㐌��K��]6����_.��k��D��|6dL��Tk[�����(�������0X�^Ć�A69��!f���/�Ҁy� ��iv�n�T�j/�+M9ض�Q��s��ϴ_�@p��
�ƥ��4�?/���7:g}.x!�����T�+b�Q�PӞ���x	���T�W4��R�T�ŃH�R�rR���C�����~#��� �~k"0�`��k-�y|*]e�?����m���O���fL��fva�
T7r`�l��(f��j�ALd�t����y2�q�Nux�f��G4D_S�Pb�)3]�A]���%H�<죨wL#�K�b$�[DS��K����l�
�dB���3��hpx.U�|>O��+��opy��9�2oUy`���� ��y��8�eu��VB�γ��v!0H���`�ڐ,-��p�M��ǳk'�r�`�cz��west?T�lc��SN��-��B��_|N�q'���(��q���>6OY����p���Tӻm W�/�2(�?BQaE�h��w�_��{�g9wA�4�O�|��z�G\t�}��I��*�S���K	V����/��������+X�
#$z_pD���{��c�K 7��~�4cn��!V�~. rB3ɰ4���*�t��)r)�d0�>����4�V�����F?�8�t}L5�5�Ɇ:�\���u���6F�n��NN���i���9 �s����8��r[¦��x[??��L���甝�k����M�l~4�KۈV����6ð�@j��agz?���b��L+��3����A�J����8l�|�S�!�"=�p��l�p��ɔUYa"je���� ��f<-�Q^]F>�,b�A���&A
�H��3I:ly1+EG��+�$�d�ݝ��k�^+x�i.������\Ǉ2�ذ�z��!�M���,���`�ؐ�`s;-�x@��ڹ=���9$�x�ܭ��M�
BJ�;���������WHd�+Yi
�C��;=^Č3/�JQ�,�턜�^�?�0���A�-b@v^}n�����,�y�����Nt[?䊃NR'����A R�����Q���A��om�)t��Og��`�G �pUn` �@s��8�m�EF�9�]��
X���Qs ��[�����A�o�"�^+�D1D����;l۵L�<�x�Y�I!4+-� E����sje�}���̉�L,�f��r�]�`�o>����4J��ǝ�v�>�p�����\Y�va�X���^�Vt���gآ�e��^+K�&��9�AF���z�-"Ys" �y:�}�� �w�i��1��
�4tV`�O�y$b�V ������$c	 Z�!r#�ﻊgh�w]\�^Li���=Rb��k�h��5���u�_�"0���)ʼ��o��P�]��z�!�A ����t����A��(H<����K�ǟ��-O8�k�v'!���Z�E{W�����ߢ�1��'�¸p&��k��4X��eX�O���	̃P���n(�ł��_�����d{�z�Ժ�7�	�N|CXJZi�Шs^���`/AI3��'�������?�
�8 �R#�Az�D��.E�K{���r�x�{�]���`�#T:�R$��BNb�0@4en�����N ��vx7b%[� ,��<�l
a r�_��o����\�Ҙd����W��W�2^H���I>��k� x�9�^h���̚�(ԝO�����"���g�Κ����;�54$4��i�d(��d���+�^ѹ�(�j�Y双-�DW-�J<�w�L�ZgS��
��qA�Z��$�r�8��̑XZ_��z���U��9z���,`B�t�'Y����_k�����W�X11���S�
yQR�]𿩘�F��^�-3Y����+�!"����9�[N��O�ښX���ԝp �9-;I�ӡ�|��~4�{�e��E�h���JTX��LP7�qvh\Qa[�,�͠�M�����f��s��p)�8+!.�ش��xO�	��I�\��������uo���@�2�5�Q-�#]�����a
��A7����_ٮ<!]��a�jIa�k��*����q�$h�P5��}_ 9�ۿ1,�7�/dj%(��z|�����,V8�[N@(��]\,�:���R�����.����+/��˩�/�s;�/�:2E��e�0��/kw�^b��ǲ{��8��"8�W�Fel���'�ȤGg�i,�n~*It��jk8{+��DD��f`N�y��)	��Nid@V⩡#Z��3�d-Ӓ9�\O���(XpӋS�����^�o�������<�.��k|?�yg�}��'�G0M�Fߍt7�)��`�m���)EQ���V��w�	�HL_i|Z���*�.	D�W��D+�U �|ԴE~���w�MF��B��p�W�$rV����ד�pI.��=/.��/�F���j�}=����3�#��D�',�3�'|�3P�����]_�O�x�Bɰ�} �{{9z¬����[`�o9��G��}��
�d��'��R��d�Xk�>boG�ATiu�.��@��Q�g��W����N?xG��{�C�hz��r2(����A\�ڷ�4<���iM*Dx]@SO�L�����y��|LM�Wj�E�{���&��\ڈ���6_����8>��I���V�T�(��t�͵�3`X��^D�g$���ො��>5��aNS��4._�둸�4_ii��N
���,����,�XA�'.B�S�'�V��������߶@�&�Ų�φ�}Y��~)/��c"�+��%�ݥ#{�mKh)�7=��M'�%���Q]Q��)�a��J�)$���u��� �H����h��%"�4k��_A��q�2�U��M�_cru�u��v��^
���ac}K�@��$�+s��iO�)P���;�Gf2�;%�����.�0��K!mRO:��fb�-�\M$�J�c(�v��J�g9A�ϭ�癱�^�{�_�>e9��dO�"�����b0�t����%�ּc��u����w��|$�<d�F'%�΃.�+��#���ڌ�1_�T�.�A��6N��"G��,M���]�&&8���hF�%^�ͩ$,n�e��[)�&^���֫Z�~����G�gN(fivH[��ȠQ\&�{Y,.�6�e]��j��>�ӞV�1�TS��"�1��V�̉��O�W��	��.G 8�ĕ�,��]���-8
�'Ԛ��;���ǥ�E��ВղF���AB�c���Z�{��iHYab3KD7"r�����
�C����(�D@������Q=��tg��N�2�`Q�3�>;�3��Af��#;�(���
�1��M��Ѽc�z����U[f�o"��tᜅ��Ix�f]���98T���1�{�qKM�2���
�6��j}X�TZ^�.�SPU��SC����k��f�^F<�Rޝ����v8���5E��ֈ!�q|FU-O��Y&X��e�*��S�-�j�ֆ!��ޔ덽�	/��"�g��wj���x����|�O��	iQe6 >ɵ��>�wT�8�n����s�+^T�&�EE�� ٧q�uҮzJ����]��+�x"��ſʪ����l�[�pc�RW���c�K\^��?L�R��y+�4=NweiR��+�4�bcd>6rN�bЕ�U8�$!���Uo.J�� �]`�9�\�+�4k�)6�W�zp2��iDt�����D� VR �AN�gqF�r�T��U�gۜ�g�"^�Ѕ��
�S����8��p"7U�z�櫚��+p��I5���r�g��)��<~��lF�m��Br2��.����^ 	LA81�2�����v��y�ߪ�/Yw��_F�� �vg�
����>�Ӟ��X�;���(E��,\x�h�!�^�O�.q9Ϧ��z�� �,O2G��KQ�W`�L��y����`��¨b��cd�����,� �Ѓ��Ew�a����ۘ]o����B��l�3?��Br��*Z��\M�W׾Ѡ^G#0�Z��bĆ�+�����:�������g���8`X��I���P�q?�\ 7 ��B"� ��&��&��{Q�k׀�P���U۱|��y����wW��0Y��ڴ�B���ۯ[V? �'����G������o[�[A��A��Ek��em���lPA��d���y�p�!�f��Π.31Z*�x�Ḕn�{]�s%�sz�t��M)�0���K��ل��r�� �v�W2$7��O��Q;���� &�I���
q��/RΑ꽛q�iՌ�Z��������r��'�78��\�o���r��V~�p.�K�3�[ ���xI��a���8�p�3u2�as���V�<�	3�<ѧ5��]0;�J@�Ym>w[��k����(���k��O�/����8GtV	G�)iOǴ�_�����=�	6OS��g�n��P�B�^B,�˻�}�ɜ�;��j;�v$2HM51,�9�6�̒q�KTb �ŔXbݮH �ƿ��g&M�	�?c�=͔��(�"����Y/9�Ť���HU��Ȓ��F�h�fu��T�
��_�Kբ��#1ٖ�;�].�ԃ��c� A(`X. ��)���ӱ���k��<�����P��
U��?+��:���	0$��TKV���ٯ�Z�̾�ѯm��7�*>�r>�� ��@̀�?�S�cO���g�������٣*����)V��n~��ž�+5���m[A4E%�$�Md)ٝ�<Ѣ�w����5��ѯ��=�@�ˊ0�C�Ds]H �)ӓiK�����Q�Z���<�ι��^n�z/Q~\�:��%�p��8�{#��f>�u�$#��W���Ij4���+�d5H��9�w�>\���������|�KgV�rf�@��AA��Fd��Q�e����ov�Q!P��$�uf�����s�u���A�j��t�<�!�a���}�=��Z��Ph�ܡ��h��\W!��X}+����# �D�ޭ�69xǋ���p�f{��y�CB��K��T��ma���'U8@CW+�P4�3&]�u�9����e&U�V�d�6��FpԖ5Ρ�v �)�U"6cZ�1�XW�[lyI�?���k2�X0��dT<>������RmN���H��aY��6�?C���}|S��QK��H��e���h�wU{b}7ߖ稵�����`�]ϻ#yl�?о��ː�D�����e~1m�VRh����9�eLpK��#ȣ����㈚c��A�g��q�����'*w.������������!eEa�X��,!�����;��O⌮�v�v˒����L�v�+��w2�toq���_��U�{��t[a�Q�/��
���uaP�3� ���Ҡ��ǆ�1��& H�
�X+\K�
@��2	�r_r7�n���p?���<�Jd�����Vlc������=Fa�q,��"��+�X�x,�P�x!�ea����a4�m����%�S� $���J�|��%.���?ͤ����6�_�׽��f��**��Ћ�P<��=�N�N�p
�8��_ѱf���l�����[�k!�WK����b`[�5_#�+1]ݲ�Af�z�X�������a('�䭥sna�Ő���{;��/⼱<�o'�ǀ׵*6�\;��"\u`����Cݙ��>&�c���`��BU"��}n�l�G@hk(��J/�F�Ñ Y$�-O�A�F@~"��������B%������"��$���`�<d��BY�s�ey!vf���K�8h�º��=.#kD)g�Y��~��@}˸��R-�P�zc~�Y@"��o<�"%�B�=%��m�[�U�?GT�Rnn��M�e���M����(Mec�:�n}V����y�����\,=��b��	ې�&���n'yY���#�]� 9O!Sp3�LB(�=)�8���~����,mw��+0 ��JIXX�L�΁����U^������k��K�獴?����ٳ���ʭ��H"⇎}
�0UJ�t��\��HO�׎h�_9��7�Z��� ��j'�}k��U�; (�'�q�j�D���rs��Ekx�!��s��.�Cl����h:��~����i�=*u5��L��)��H��-rV_�'p�H��`��/tKmBn�?M1�C�Z�6e�2��Ҫ<_�,Rs9�g����ե�8.�Ssg�"�4�;zKo����cAS�W`=����L�W��o8֟�K:��I��	}l\~ LA`��s�Ԧ?ۮ��BI�y�5����NT���\��h����o���,)<���r����S���x���{�|�4��p�{�?��{��j�\���cU.\�Qs����'��`� �́�ҩ��]����[�^�SQ����ﾲZ��ìXĦR%W��NI�C��=-`�������<D�j��تL����Ҕ����):Y��'%Q�*l�
�3pE�UmOK��>E���=7����;���qt{�����2��B'�}��wc�����k����%"Es�@��V%�F��3~�:�-ھ߅�Wi�!� Z��!�(۪��A���^'����!O���4���>o	$ٵ)��L���C�GbXp�x�rݰ@���2�ݩ=.�3�/v�J�ݑ�Nc?�'����I
VU]��ث�f���Gg�O>~�2���lr<�AG0�б�>��ˠ����R�,���*�;�mˆ}=*�B���bJo�T'�g�c�����r��dLڛOZͯ�¼�S&]��)���\؉��L�<��B.��'�^J��:,�ך��9�-Т��Ģ�������Z~AKg�'�~��F�c��2(Z Q,>�I{Q�葜�1��"�#�2 �I;R��'�}4̬��z���~�U�i�$��ݸwBe��~�[�SxU��'��l:�,|�q���[�zug�5w\��Ԝ�o��K��4�2�Ԅ�]6hX����6t7��G���-��]n��U�n�r�ñ��>@��iɛXp�Q?�A����j��I�S]�~��m�<�s^��Q�]��X�ض/��Z]zڿ����mG���~�E��I�>�������������TqY�Q�g��ц P�T�d��5Qq�+�-�/�J48��PF�^�����𲆣�n\B 2���5�M�	���gg����b��.��3ԠQ�6|��m�Ŀ����w��f�0��٢�9�ԍrƑH��P����`�a�"�p ���J#"��ۖ7�g��U�#�δ)zY�����`pvx��V4�?�A�O�|�`�
������\ �|�}4�Q��%���Q,�xV>�����>�����T��!�fO$�L�*~HD���L���q�͉*����n�x���"S6|�]���6a �z6ߙ?)z�ʏ��Q��Z�E�]��B�����udr̷u�(���?�d�J{x�cA����.����P��B#�A1'*_��5gp���W>��QP��Jy�� ���0�r�*��5x����x!%|�NZ��=W�6�o-����#�]nb���)�Z��`��ܿ"@��c��s�q�����~L�]uU5���VE kR��,aj��vsp��%ls<��ӧUj<8޵�nQ��SЂ �V�!�VȻ:4��/%#G�d!��y_��3����0�7�;e����lX�dBɀZ�S0�nuBZi��C����1��|�=�tuN>�p9*j���f��a�bn��j�цW�{�o��,>y��F�es7{j�j�|ܟ�1د� �� ��52�w4C�TW%��NJ�4S3�0��$�=��Ǎu��oM*ٌ�B�_PK�������WH��.4�K.�ߝd��� } [M@S�=?<+$���5tg2(>�|{�e�Y��wL���=�ᆎ&=܊
�9��z�e�;U����Z�EN�<��[��B��|���u<�S���}���v�,�<]:�qHhh��@U���O���$[�ϕ����f�#�>s'��CK�)����,+�����h۟���v'v	��3k�(��Q�Z�H��k�a'�Uy�ps��d\w�D�2�N��	@S0��B<(��F�Zou'�3�<�>EmH�8A��%��4�mgl�8k��s��xN ���~T�-�ZS�r.�z{�^���\\-$Ն�D�ʹ�C�\0uX����h��Ѓt�Yֆ�Y�l��#Za��%<�}���]�}Ť�aQ�^���x �p��Z�m�e���>���ȑ
�������I�;71>l�0$|T(�Q�ֺ����|cg�2᧑~����A��[�>4l«0� �0D��1U̠L����#Y?�:��*�I��q��T�Z�<LV<4O6��w��z�����6BTĶ[��$���2����I c����^l1{����]������
M:���B���4)FE����W�~'�C��$������V��/�W�3L�-�0�S���_�l �]�O����H�h���!u7�~R?���*�r���x(#
�0l��!�Њ�~�.xJpq:G������w�%@�_�1��`^U^�$�?!g/)F�X �t%�@��p�7
(�O7�,
>)��Lq�B��2��XW��eaZ�� O�o2}<�0�"(ͣ�� ��ä�
H�՚�V��T���F776����CB���Z����Y_M��k؉���]2���d_�\Yo�VN�_puY{@������ ��?G��F~d=���� :��S*I�=;TIwŦ�����\�ܰ�69�,�Jg��V�$K��TeL�>����1�7Pם��SR�1�l�;��������E���;*�%��^[|�}���O?H��Q�.�x�8�8�HJ�I����I:J�1��V,P�¨'� �q�/��.���Ns%璟/�Cl��<�S�.D`�]yY�kAZ�qd/��6��$�&xGc�S�#Z�5)�:^�mU��f� h`��&�|#��n�����5���piQu� >�����ȧ���woP��朁�DV�A7_���t<���%͗�7Rkݣ&�D/���!�Nݟ�3s)#-��z����K�EEXLz�XZS�t^�Ak�+�n�����w�1��	�LF_�+��$�g�[< �m�>'���������C��ƌ�s�X����A��h��"E�T��{L~B j&(�=�g�	; {�Xu��z���k<��9U}`�� �o�z��Ŝ��oJ�SD�&����2C�n�%?��F%W�5����xf��lŘx8�7��"Pz(�x7�?W��P�������<-Vg1� b���#���o$���/����o]�g��d31罓�������9I���8[Zˌ�w�ϖ���m��R��0�y��$(�~�n��c�mR[�X����T(�Ӎ�D��}
{
X��,S���_��.;�(�u,4o�W,x��.t��R�x���t��A�&�Z�Rb4V;��<J���o�=�$�OS��A��u���i��}:�/䂴�f74 OTc�h˺��L9�5�$��~�;R3�Hl@�B�J������MV��P��!�*C�{���i\��7C����E���ؠZg�-��"0�I2˿"���w�V#�зg���gC������'�����w�aI�^�T�Q*m���6�F��Lo����"�~�]y"��a���I��x�6Z\A�+l�$5{%N��e�w�kX�7��@�
��~Oq�z�)F;k�����j@q���7	,ܸ�짶���_GzA������)ԧ1]��t�ڽ�7A�+"�V����i���Mf�(Q\�Uo$��Z�������?��|"��w����f*��fD��uՐ�m%Ue7n�����.=�J�m��k����	������ڕ�v�<'�d2XU��r�x����"߆o���À����U��Aj_,}�����\ݍݹ�n�*�t5���/۴݂��H�M�_�m�L�Ȯ�xy�k��yh���ڔW�� �s�$\}\�v��O��S��4[���3m�<nܩ0?�o�%qU�e`/Yw��=Ig�a��^@zL*n�|��0K 8+�MJEE~�#UT����t�m���(��/E�>*��}:�+�?�9���P�"��S�:�3��k����tGG�%>��#d���֔��IJc��W
V 
߾95����A	ݫP�W����
TW�X"ٶ�y}��Z�� $.!@��(
3(���3%�j�@�d�h(!h�?���B=Q葞�Tߚj��O�L2�6^���T��p�^T�n^f��\7�<3{�B��Vy) ����l�S�.U�9ڸ�#�L���{��P��n�`}�e)��y���4��ċՋ��%��h�vП:`(��H�}�;Ȭ���nS /�E��k��&LR"�3����&�ײU�*�Uz>�O���1��i�h��a/���&~�����s�|u�kC88�]�xW�3Q��JTcwM���@�{������@�;������(�����I�A����eq��n��,^qm���p�23ʈ:O9b�6���K:�G?�u��^�0+n�]ʾ���]�2t���{ߥ5�"R�ǛQ����W=�t�Q�0����i��O�0��
ߖf���y��$�;�%�. �.=Ч ��QG}vc"�C$�#�|�>�u`"���\�w�3���v�p����ȵ�R� ӼYrf�%e�t�X�O�|g�a`���h��c&P�u�P=Vܸ��_u.��4u�C�Zh�i�.j|%M6c2���L�/g�J����͖��9V�'��[Ы�_�{LhۅD �q�3��V�AoNz��"���Eى�Vz��$(k����9�j�Ւƅ/j�G)xЌ��-��:U،�$nکJ��7Q���͏��z�o͊���p�s�_ �$�0��{I���s��T��?��l`��R�lڱ�C��ٕ�QK��TȇNR��0�|�.�";�2�I�d��L��רh,�L���p��L �)c=��� ��]i�nc`  �Zl��{/�3��dɏy�S[���t�M�AH�X����|��n*K�C�2�y�d�m�T�����Ħ�˨�)d�~/_�)
������E�-r*�ĩW�]y�g��N	��|�+RP����?T��]� ۨwEtz��E�%�uµzLnӃ���@��b�~�'ړ�T�� �UqDv</�F�J$�\�>I߬���S3�y������
K��Dv�B?
\�H�󆺞�*(��U��ߟ�i���$�^�v~��ހN�.u�i}��%Zv�ғr
;��HB�0W����$L�H��Lj�g�N�m+��@*��񇴹�:�*���%*��d�Ȋj�5*��!����{A����m�d�;���QIN�N�P=�^�Z�"P?� �za>lK �0,��t����z�����r�̸xڗ�j���dq��e\�­�r�'QK}�N�]C�
��K����l�n8��
V�y:�wƀuTɝ�&c�b˿j@�)L�d�@�+:�a|�.�adE�����$3�7�^+���]�޻&cNb�ժ�4a�A���H�Y�wl����q�m�\��-�Oў\���}g�׿�UtB�)[#���t�#
r}f�AD�'ꢇ�\|^tz
���=C��m"��"��ŀBGK�pb��D��Ӕ��=�j˷$��r��&��5��;��d���Z�
� ���;v��Ҭ�R�1'�~oQ� QP���Uܜ9��e#
��圹��b�|4�`KNZ�䌴�MŇ�S�|Oi4���,׭~���C���ys�DU��۾l���t2�ǶbBY\ܨ��moO)`�C++!����	A�ݏَEb6W,㭉"�e�݅�7�P��?� O�l�رZkP�P�R�w@�&Y�rw�h@�V{qa��N;v��j ҹ��������0�Ĩh�iՖ~��[�.�
��V�c(��)]x?S+'�
���w�ux�^-��">z~��B0��㈫�V�/e��F�Q�[����O1Np�S�{��H#�`3���3�uz8�0�X��u���6##De�͸Ƣ�yg~�J,����ʜe6k�������.��n@A>Ȩi0�y�4�[I��
�aJ�S5"X�<���t|�����fKġO˲��{4��N�Ʊ��
�Yb�Fg}�SB�s�р:z�g���C�OGq���̡qt��4R $&A
v�\�3&\8��5�UT:���6N�R� ;G��~	�r@�匉�d7�vJ�#h�h`5�&���P���A!�i���/y[,M�c����ϋm��ս�
�(5��qM��N�IC�@����;��nT6�α��E�;1�z��A^	.V$	����@����N�aDM��jm+g��)Ƚ���jd6\������J"�Uj�n��̿�e��SF�i��=>m�H���ٿ5#�n�k!����@-:,)��.E�:B�%tgv�ի�)�X �TP���)|�S�
��EY���~��O,7�S)��SE�?,����*�,���DQ2\2,..ZQ��]>�8��`[R�`�m��z":��{ی�B
��\��S�\S��[��T�������ŝ����.�ҍ2j�(6�Ⲡ$���ޑ�_�H!�a(x�-�p����.��Fld�0@��O=3Iě`�ȌbԂ��s�B~���D5�nZ�F��ëL,T����EM��7�"tu��\	e�H����+�Q�YևcX��2����.�JY8���Ç0G`�"�:S��[�Y��u���:��u�O��򁺷4 -�G5���Z/�Ov����~'�X��%2h�gj��6�Н2��?���A!v��mUj�ؔ�UBBijk����Q\}�K?�a����ŝ@t�6�bg l.�ǐ�`�2Y.!��k��+�^��8����q��(Ͱu�k/�	E��������b4]��[����;ё��K<�4z@w��l���\���#�'�G�r�^����;���;��>*Ћ�!ߪ{&�>T+Hµ���d��2���>�~E�C�ߴ��&j�[J�֖�z��V��Y��f�ቓ���X����?���3�	G*p����؛-x�=qy���<4�wD��X��uՖl���v
����&�	����+p�\��
K�&w|Cn��`��G���%�R�U���+���L����?�B:��!��h��g�[!$�p�&�D�#�J�"&`D���O���g��~Q��{)S�YnB	N^b�ݖ�?�E�h�3���mQ �x��"�I����\P���WGdZ	�oSe f��̘݉��`�*�SA�Q��6�Q��噙v���\�
��^��x\ m���|$U�j"�c�&���/w��D$���ҋ�8�|`~_�v���]��8�#�����	}�]��ӏ�Ip�3Z�?9�@�^��Ye}�+���kIb�H�ւ�MR-��j��pꉤ��K,�ٙ����;�s2���� �l�)�>	�;-lL�(��,���E��d�:�\d���N9r���QM]<�I����J����L�x�P7g�
� ���'��hvL�Ѭ���D�Saz�����דl�]��2s�t�	?�`;5H���9�%Ѱ�]�v�ǈ��sF���!�xq6�V��ݚؒ�P7k�Ee@��Xu�p�8�92���ۛ-��Y?�JfyZã�u��,�)�㑎�Փ5����k��Ԝ����2�2���n�08ɘl�����N�6��^��#z�
���.	E8����K��W�5\; vl\�[�!�f�>�='�ջ#�۱�uW5$�}�*Dؑ�X�po�,O�K�Y~Cl��m3��y^1�\N�������Zߖ�PB�EYyZ���-�2��X�;��5g�0�GI�u?�%n��槖i��a6��E��6n
��$fb�S2���l�"�U?T�W�`�~��e��y��2L��t�,h70%D���X^=5�4>-��"Q��ĭ�OF�?�۽�B������<7^�3��Λ�HQ�ɇz4	�&����Kk����(f󥈑h��PL���{��t�b�q$r#�����C��S��Wk42�N υ�Lۢ�z�Г<*Q�e�ӜP%&�=`��&>=��hY*f�I�J����\�[�޺ؤ^DW5��y���v`ܸ�#�ҷ76s�)�r(��X|GTġ�&mx�v�H��)����:D4fp0�h��������b�Ekw���Y���!�NY�HN@�U��܏Kq��*�J؋	|����}��0�������T���'T�����k�,���{��vs3R#���m�n�cnk���dd{��G@�"��L����R�&���Ӡ�,ߪ8R��M�H��[	�B	v���ȾO0ɿ�u�W�5�=�����D�������N����>�͙C$�ɜ~�f)H��_v���x�ޗ"_�c|�?PL������Z���)kZ�����:F
$���z���Y(���������/H}�C��܅=�\K�	��� �t�}�������
cf��Ηpj*\�8oy�C%��CѢO{aFġ��'�{��vp�y��C���u�I�� ����2�Z
��J�x
n�SN_$��A�S��\�8d��4Lkݔ�B��2��n�D*p��4�S0���1�~����M���/_#ţ�2ﴴ�9�X��6�Ճ��ۂ�m>d������o��9�w!�hڑ[D~���HM�����c�C\��K�2�1�]�A������r��	���J�Z|*z�4�iF��Y��\S�|ޘ�'"I���>�93���ᑺ���߮;3p:���K ����!*>�>�I�í/�l����W��q��c������i�s��0C!��z�y���T��=<.��Ǹ髠�9:3��X��[��
��&��Q
�!Ns��}�F�k%��� ���DAvx@���޴WX؍|zDWϙ���h�������_|���g�mF=�t?t���V�,�d�$�wUc�c"�$wY �((�͒l_ۣ���4�N⹟m�MC8S���G�e���q�$����֧���"E�����j�ǝ�/�1tn���<�GN�rT�`��Iz�X#������Hlet0o���~����Q{���R@2 ����6oRN�+�q��5�Wk��4.�aH�A�ph�#�7��tv�Rz#���Η%N/������2�����dsrZ�b'��&s�엪�0�$>�C� ���k�H��ۙ� Ȱ��
kGf��I㫕r��sDo�jvi��+n5_���Q�B��I�n���$� 0��:G�<�Z"g��&ƞ�Q����{������T<8!��\yY�X�-e/��7b=)��@���[�o��$�E�[K���&�wn�"��|+��]�j����3��6Sg@������_რC(��BD.��NZ��T�n�>@֢	���oé��rz�+u�oʭaYwi��hd��ˌ�����*���
$o�K9ל0{��r`!��i�0��]�l߸�v%8o��$�ϊ���F-���-U��8��,v���ߜ��2��IY�G��ujyL#���ҽ��⬙���-TS�<Jdm�tp��\�}�gK�Y���&{�����_|��E��qdB��+=����T�Z<B���I!S�+Y��Q�0z��e�
��=&?���`�߫3g��F��o�5PA�6��������bΗq���"��ʫ:./�P�L�/�x���  2�
�\lf��\P��:����Q^I�-�k��Ny�ܫ�W����v;'G��fbʟ�F�ɟ
��T
%�3��`�{�O����-���oކ��O�o%��k��f��
����Vq�\�|��o�Y��F[8������56��/���l��KG��#$ �m1�wJ�Q��l�5�r!�;!�P(�AU&zͲS+
\��!�k�6_�ߨ$�N9�W�8��D���JtZǍ� ��|-��٨�'�Jb��S�"�T(ۇ!�,�Cp/�����:N�f�����}.�P�^��uP;��������>�2W�H�Jcf���)�O��]���W�1���2x�xdM&�>�4g�x���~��'b�b�Z��c��Ɲ��m�)�?+���#��+����1�Ay� �*8X��"Z��c�������y8D9�S��&�o��7Z�&�@pk��^�<F�r3\�m��7�UW���5�,R/�v-j!�⠳a�3s�r�ld;�3���˽4B��O.�#��$i�_�j��̐�w�ݦ;��:a�n7�,��8k��~�>Z��ހF�,�=.e�V�>����I�9��J���)���=i�D�
�a�m���Q��3wc�N��t:Q��Lۋڦ���7�S���ȱ,W��ox�I�N�� ?Fh7.���NzBKn"����_m���s'�.줟ۃ��J���*$���y(�Kd+}���a��+g�u��b��=�K�Pו��X:�L�+H�7�8��1����i�8@4��4�����ۚ�j%�с�JQ�"8u��:=�e�sz斋��W�r����L������>U冢7il݆=��έ�q��C��t�{]�FSr�/�{gE8d/�_	{� �f�C�����@I��}�@����߳�S~�'ʠ�O�gZ�͘2�!XgO���s�	�H��F��j��H�y`�G	�Y��0A�2B�_r���ݙ�V�}��մ�d����4�x�G�S��|x��P�ӄb�O+�L���Ē�}9�Vg��ts�^�U���_g�3�&�ġ� >�(�ػ���/W&�Ƅ��U�z����`��|T��R��^���΢6G�s��ıl���s���p�*��h����S݉��ƫ/��tgG�V��y��FC�VPmv���3R�L+s,�$P--="�)�5��х�m	��<���y��M����L֗P���4��Y�}�d����9���Sp'B8e4��v�� ��]���cD��;q��.y�+45Y��A}&�`��~̅�}�[E�5o�"q�����))j�^�̓]���/��5U����	-	��_}�!=���BA�-��@[CM���B�]b�
W�O��H'����/$�N�Wƅ~��a�5L��⭆�0�$��޳��*�OR*'v��́�>I�l����u�3���rq�y�-Q�ͤ��3�v��s%t�1&���ޭ3�7|:��������uG0���w��9��Dg�m��$O�~���!CРX�st\��	�����'4�O0�S�\t��QT�`#��L9d�{i@��Ĉ1����Ay���}Ӂۛ���*�L�6� 6�\ǳ4��Bn�J��o�_k ����WYb4���@��DsY�;��]�?࿖v� ��k��c��c�1c���3���P�n$_b�#tΌ^�@��""�Z�eGq?+�^xq�v|��}Fj�|Ky�p��qM�%�P���U&�rV"
M��w��q{γW�z�L������� ����ډ�#+�P���$!:
?Ca=`�0�kU�l��䬜N�Ly��}�t)�������l�Q-���?X�Cj����A��v�fsI���e=��JN�9o�	C����)�FL�nm��0#%���?P��M���8�Y�%G�U�³�����]��Q�����C]��<6�LI���PU��w,����/��랶�S�y�rM��"���n9��N�\�wЛ������t������x!E	�m�� 1��FG.4�	�=��8gk��˻c&���/�X3�d�541W)��w��,�/׉�HS �9x[1lߑ��a� X}�gU���ꖡ�.L����W�m-�x}���v�<�����8h\cyd&{]����rYwlέ�8!8�PL46u)�Z��<�,1�4�,�j�j����VwuPg����GU/B`I<V�V�_�1�̀��=�й��u,y�A�Ur;+����B�eAVWC*P��V����Ȉ���b��x�x{����V�f�JJG�?|LZ�=��d��ȣt\ZJ�-�I���*��T�����O��]V^6��$a��$b\���\��$��E~��Z���a4��v�0�F�-�0��$�O����UV��U+�*�G
4cg��`��.�� rԽ�e��b��kS����N�D��&�A�"�eU�c�+���^�/�]�6U��?��6�w��I��z8o�鈜k��%w��(�:JPWۗj���\y($�P�8K{=���^�I}�&�/�f^F�G�S}�`�3������S&"�����&y ��WT�A=����b�ѻ(}�+�Y �Z+�������[�t��|J+�U�{��_< �>
�G�V8��M�,P`o�vu�c 
�'��#�}Rj�G��U�`5X��L;L���uG�'���� �T�	S���)JC�,	��5��]jmC��, ;�������,����B���Jj�ږ$�!��
"�G�q@ٺ�G]���q[��!N"BE��ŀ:3$nf���@��˘�h�+��ۮ'$�LYP*@�F�t�Ð:c���ǐ	���4�!8<[ڵ��E�/�G9K������Vv ��]���4����J�����̷!�,�x�v�P�|Y��fO�0W7*�z��on!x�(��C$�aE�R�
78i�Rˉ�X~���ҭ�K��J���C��{�3D?���R8M���8�#�T�F=`JEm���[@D�#�[i�%��]�H:$Q�D9�)4l�����Hu������G�Ǒ���-�_X�w�T�¡A뤦v�����@p��W����$(��
忙/��x�plp���s�w���῟-:�\�8b��S�?脄�?�:E�*�P<��Q��;����Ṣ��S�>@��>�����a�Ck1�
:�aZ�rL�~�w�ۼ$�$�걠�"c�+R��f�wRjʿ���i��f�ƻ:II\N���r�/�W<Oli瞫�x�<F$ﾩm���'�F�O�.d��9}���Hf�^	���:|���UԹ�mY�k�"d�������4o�l��ި�Rb���l?8�}|z-B|���ܣ���'	��K�D�J���)v��jO��wWmS,#�X"i�)I�4�L�Ɏ%ɇ�b�l�~E�������g:w�U�g+�<$L �N��l�їHRc��'�d�W������_��~8e�$⼗<�)\]du����F�H{�kX�x�!;9י�tr5�9� R/�Jh�����E��thS� �ǆj�#��  jͱ�U{�Ll1#�y��F��}'�hs�(���ꔒ��I8!5$*�A����+�z*�p����F�%�%�z6;6Ĩ(8݇�.(^%�*eܑHt���_�x��5�c�g�Lc��c��[/(��b�=����M�ޔaè�
��
�O��_��>��u�Y։̇�h�=��l�j�gI�����]�M��N��D�A��H��YY. �W:&�j�u��4�����vxd;�D���FR�l�	����G�Kx?�v�g�Dڪ�;�.����,�iZͣ������h�Q��/��.z;֗b{U���}Rܮo�A�G8I����i�F�,��n���q��=ǽ}x���k�Hd��?Дї̮��Į+�׌���[K�c�����*ӧ�15�<�k�����㹾�A�ϱ��fʀ(i��uz�H�fj�CA�P�� xp
�>+1��k�]s�r �� 5%hSC}9!P���;;/�w�����m:]�r
�7��㼫�.���U�2&ZKo�j����
�]L���������ݺ�Bg<[Oޣ���!�U�ݶN�v\[SS�i�YjP�^!}�)�N|��}?��s/�tKiJlx����8��/���UY}�2B^�<W:����$��P��?L��z�s����<�x����ޢ{���Pҍb��II�s%J�,�c�K�]q�ʀ�)P-8tW�����mxNCZ۞�N+�BQ,f���Eڌ���f����࢔F�(5��\���>jh���d�g���fh֘�g�Q�����ڪ���"	���h�\'5��[>��DS(���*%f�Vfa�d�8����\鋧nbM�3���
sl����y����WZ�n;�g��h�-eryk=ΰL?�w
g��7<�ƥ���x��}�ձe��+-����>pr/���?�h�%ݰ�55d5�1�p�"
�إaZ\ږ"�^��ϩI���/�d8��$�:����a;+'a$t��FǾ�YE��S�\���_�O�M������ZDm��B�?&q���ӱSu�9�k�ܮ5���(�i��SY,$9���/�yP2�]�'�n!�$��J
�f}�f!����0�n��/{CWP^^��|��������M��z���$�b&�wAyWw�)/<]�kW�+�1�a)��8'���C+�R��!e{
���i��0|�������qB�ŗ0�H�2�\ڣɫ�<,��ʵ-/m�����$����	�q�Y��UQ�?6�z8�o^���L_���&�]�]B1D��-P/��g�.�n'N������_��ES� U*.�A�u����a��)��_�7/I�>?��ډ.�GP�`+Ν���pM r��Kh�|�~77�}�ZH�����^#���o� �C��7 �,���`��j�ݵ�@9��<ܾ��Z�1�~��Xv��>���z��}��X���3�7�'e���:;�&���/G^��T��]q���7�SH�[�4� >u~��Xc/Q�;���3A�]qO�[b��vmH�H�uO���� ������p�ϵ�^ ��X���U�^ ��
EG��GC]{�
u/�U��h�ڨ���*�dcg@04���a+T�Drʏ���@y7�x˟����Q�9�������g�o�P�?�0
��Y�N�\�+��m�B��o��/C/�����*� �:|op���x1�gn��oBcT-�U�z�k��_�Z�Ҟ��C^�&�#�}s'�N�^�:F �?:8�:� jKM����u�y��{�8��4���^�:e~ϱ��Tt�0���ο���_��t�jƮ�_c:xsdJ;o\0�|
���&Zu�����*�-���Jo���M>���Ĵ��FI�*��41Rl��uX�e�E5?slc�ZNF�[Ҝhq���U�\�rt;FaY����hK����׃X�[�ڡEt��M
d~�=�]�.��Y�NIg�_�T�[;!����b��VҎa�o=�s�)��v�$�6����s��՟"..���Hc����}���7�}�R��W�3s�t�ķ�[������,�5�	ԁ�Tɛ�OC�����N���|=�.��3yy	���aj����7e �Eaw�ck��b���;zBYƗK�b��e\��UI{9I�/��7�R��
��,��IK#�t��mOZNl�?��8�̾��+���e�3-�����D�ٳM��O����Z$��|�1ic�POທL��G�z]M�����������q=�fj��_H��9���>�.| ��q;����,�3e�-����j�?���#�r���6)>l5���������J�\�o����P8:B��zmQ��Sf�)ٶ�t-j�P 4��'i�<��p�J(W��vCRJ� S~Q���g׳q�wu�
ڔ�0k�F�����]Dw�686�ydu��[w��D #"�0[�rC�	
m�D={;�qS]�͎���,��0��T+�����|>ʛ�] q�F�@���R��Pk���5�rއ�#���=����9�g�������e)� X���6�ӥz�X�������z'�4ʮy��kOG��+=��O�s�8��D��M;�P�U�	�QE
��0��OY���{ᔧ��{=����(˗���ތ<�B����3� em�|��>2#���1le<¡^��̅���O�^H�}���x��OeHá���¦{�N�|�H��=x��4V��چ��vV�T�$��?H�`sU���Y�@���g��\X��=EWd��}������&�fg�/�.uE�\j����u��A�R�.9��[!OK�trF��$pl��@9�Z�	�s�~j��qG6�uA�	"]Ga���6��X8n���̽�Q�.�j���$h�g}P#�;`4C`�� �Z�����n��u"�y���|qZ{1�m=eh��	�}H�z�^6zJ/�I�����Z6%cy �?&y�̀�S7=1���֩���Ë�RM'���?q���9�X1����F	��(��ĝ�e��L��򬹵9�R��-�`]z{�簇�$�b����Ng�(w��قr�m��I�|�,�&�˔��DK�<����������Vo'�{)MU�u���lsߎ������zk_2��i���-`�p2��.:.�����׀W�?�I���������_}m)!2j��L��{����Z�Y��~�����S��:�E��`���𻬨!��c��}R�w[���.���߳�?���~�s���P@�,:Bn��xY������`�C0�ab����}b���n�����mj���M`��ۼQ.�;�.�1����m��w1U�'2�Oq��W�9nD �/7ɊYW�����êL-���L�w�dbC��lS�7�b��a"��C�U�@F���LU��^�<���!�3?�����$G��m%>�m�Չ6�VVe��rq��G���a	�Gx��n�J�B<��Z�l�?a3�e��X��e-ɒҐ5Q~�W6g��WY(�s{5�R�H�	��c���A�/~# Fc�HZ�: ����4�}�FpHmR�hU���BR��@��kTf�z��do^�C�֦|���^���_��N$o���l�1��V����7�`�������͐���7������$����T�k8�
�Ϫ �T3�G�B��#��6p@���M����g 1�v����h���\��FO�哽�'i�^P�_&�PIpGZ�ta�#�3�O�]�b�y��1��d��v���%���Nyc\+�
hݭw�/�c��(@0j~�����n�3���)�4��y_�[ v�����L���A<��5�GB2W��elTa*|����2�<(�-\+���ӡ�Zf0۝f^6"����6G;f'�kR��N/�g@kܣ�.�I�����#��q^,p�� �E�7}`��l$^�ϱ3���x���A]@)��A��ѳ�
o��诇�����D~�W�z�I��az��?G���
GdA�״�<e_�ТC��*��Gx(�ƛ�B{[����Y���Β�����4�tV��å�G�Rͯrk_�Ӏ���-����~�ҁ��tP���w�m4 ����w�e���&E��@�L
DQ���Oφթ9�s��q��e�Oܜ)[�P˫`�z=����=M�ft��0�x��UTˢ��P!� �2M�n�%1�0Ŷ�|/SY����b���˕V
	����.���lB�-���#���8�{��Ab�N�L`	T�#'P�E'�V�I��;~i�_D���Z ���}�fN}���9����d��vxf02�2��|?�]NV�������,���[�A�أӚbV�r��չ�֫H�>7�?��-�w�o�m��r׫l��~�pZ��~�+$y�]��M�w�ǥ���;�ۉ��O�R��q茄�jdz��wn�#QZ��FP����m�y����v�_�[.4�6U<o�0�g>fA��%�;�9�V�*c@�����r���p��P��&R٦G��i�]�#b1��>� �7����q�xɣ��^v���S��y�.ga�������ߑ ����ڍ��)|�R��'i�|5Ѽ�gAtr�E��4�����Ztn�q#J���,��e�S�	6\`%s�����:���F�����*���L���f��>nr;�")[`IY3V��5�o����avj�Ƀ��P�T`�� O��/��'�f.#�pn��F�j/\5V^]f�?���7�5)yiG������7�}�)V���5n���m/ �5���#�x\�-j��Y#6iJ�(F����E�=c���<3��'6� ��088������I%*�i� +�����~>����"s�_2�d���2O�b�h���d���j�r���HFW�Mp�h�n7fRrf:2U\ uVAЦ��9b�K�̽^t�Z�:�yW�	��r�_�:q
�x*�8�Mu̎�:��U�{�;_=�D�h&� x-�UjΦ�R��Eg��	�b�-�������.ZbO����S�^�uNz�a�!u�����2�4�{��A&�e�7������;��x(U�6���`�~!�o������#���/t�Jr��i6^�W�+:<R-�o�S�> G����VxHB�������`-5a�?�4m�A�����UG5{^}xځ��R�EQ��m���cc�c��0�ۋ��{���@�1|���� А�%���z�w���X��:(?B���@��S�Q:�����7��\��"�<�}��0F~�=��-CZ��j�F&8!@�QA`��8��+ТǼ�
.w���C|���� �uiӛ��l7�\�D��<<GD�o����T�~gb8� VF %閁f�o��0�hP�T.���v#��gJ��,��C��M��
b>�P ��lg�z��A�T�`���66�{�}k��<���-	��0�c�}P�.���I��Έpx���N� ;�,"x�A�Y�Ӷ΂ʺ����1��{ޡ��d�Ϲ�8+Oc����I��G��~�-�	d�c��J\Q�$^��w�+
����dxX�VwX&�#CX�Fh:pP�;U�5	+^F���]������?�[��?���! ��%nh
a;����2��J�Q����g�]�m�^ �V#�ɍLmY�Qҝ�F_D��N�J����;C�IgMn��GKܹ6)̈���:�^�(|6��<�%W��h��rׯ˨\�˶��ͷ�D�����������©�6T�V��zV4���}�
9sLF���O|l���^�$r�Lf�U@�<	i���l���Q�%��卪�s��~$�V����~�SYl��Υ���X�����	r��&�'��]*��)oe�&+{����|`g�beY��9){��t1�ݏ]��ۧ4��c[T�v'>X�"�'�g�2d�l�뭛�J�]7��X��+�W����:��u�!��|+�)6�X�k��vsUQ3�f��m���ǅ�4:J�d�hצ+�稭��w��'�{(~e���#�뷳�_r��6>�A5���Щ4C���H|�v�.<����K��Ԙ����v�
�fk��{9�}m��X����(P:���;۞P^�7j���&|�k�cЊ`��A�[`J{��{�S'f5�&�	l���
u����
�t���k|��ѝR��U��V��`k�ܽ��@U�Ő|n��n����	��i;1���e��<)�b����n�X�&�p�62��ޱq�reNS�iK8��d��ރ��VVB�a�b	b�t��/"�5y݋�^�f�.hux���3w�/� B6�R��Of����U'nʾ�����XLj�>�� <D3��r��tf5s[���/Į�8�����ڦ�Y����=�w��@�tH2�n�]ߘ��<���c�~��e�c�4+\�����\d� w&�����E��Bq�o�.�O��8��?�iϑ�0���px y��R��iDh����dz6�><ߢj���cM��C����!K�X��}�N��-���,�6š|:��<#=T��M��x��$_"M(	�A��P#�.��*�x���$������\�d!ĕIo����`m�Od�@)F�яIǜ[DW`*E�F$+Ta�����z��[�Q$g�(�ĉ��eUS����q��Be��6j�hvy#���m
��c�<�`a���.��u��i�"n-܊�Fl�����E�ol��j��8[�Dm�z�-�è�Uq��t����T��R��.��I{�o�|nW��X��qL�bG;�cl�Xҙ��� �����;j��}�j�ԕ��ܔR89��k�m-N�Z%��B�
�A����d^3�s�,�W�����UA� �K6�o�,+;&ь룖��s��E0fF�i����0}W�8Z ����WPW�e"�hN��ٴ꓊��N��lu,]���P��vَ��Y4����u�o�4����)��)F�6�y>M�Ef{�J�1�c��� ��g�\�nh�	Ee���Ѧ��e���0�w�w�Đ�n��g<U|�# ����"8-6o% �)�pF	�C���(�p�7�a��{pֱ):��� �KU���_ ���颩�;=%��6��.e�� �8�4їY���v��t��4:��L�˼��?�F��|i��B���8(�R�@O7E�6?&N��f`  4���li��>��n, ��nQ6=	c�#���?�u����E�X���*�S�	5�!�M{�GL�P�a
�����{�	��b�_���݆W>4��[Ο���P��mX5�q� `��P�[y��F�+�Dc̑S�/�'�e��e�t�y��Y|�7�TYG���.�1y�oZ("+SeA�R�.�DX�.�7b4Oj��D��b� zj�����`�Gg)�E���Vd|ڤ�|԰$Q&�P|�0�*��2G�LĜ����+=j��wMj�1�E9�*������W������Iv@M�ۂ�ۘ�V��D�s6�^�'���K#��g�v� �r�'�xi��b��.�H�R��W��s��2Y�e�LN�5�|�n�ӻ� ~��̭7���%�'�T��I/m�c�䐅�Ј"�PQ@��f��h�Dś��gl�LS�˘���1�Aq�P�f A�C}e������.����ɑ�	���l!�Z���zʃ�����_�>*O~�t�[����M���M�S016��2�@�7Ɂ������p��������v�y��j6��Z�b5����}��Ԉ��h|'����T�B&�����t���0��(��[2�Ȃ}����0f�K�0��|�8��r
y4m�]�Z�X�u&�L6��Ưp��KޛٰqŞ�׿Q��!���|�����U��r|�T�Zo�`KY��,Ģ����Ϫ�k���iOB6�IW�T{��t�:��w�ygyZ�������>7��0�$�qK��,�?2B(��넞�ňGQV^1�fЫ�IUm���S�r�ǆʍ1�� �>��m��� R����c�$sB�.�`Ɠi����:a|Qb�O ���Ŧ�����A�v`�P���\�NI:]r�ы��L,����lE��H��N�Cޟ�Mz���7�߻C'��m�
��o	x9#����4�Y���4�JI�>�uT�#��3}�����p�L��k}/آ�A�wɅw+�W�4A�[�g�^?9�wi	P��_lW��Z��4�b�)�����~B�帯����\rJǎ�z	#i�%4�p5.\[�eY>�p�a,���ԈE5wS+�D@FX4�����qdy7���GiF$�l�8�g���9�v�]�F��hH��[8Nڸ�������RZv���1��֣B�Mr���/ɇV6���j@�ǃ�T ��u!|�K����~��N��#	���c�oŧ��� 쑫��;��{�6��#>�8�Н�(k��C�J��Ӯ_�z6�#[�|�@\e]���l�#�c����nK ��'0B�
gי�-�"t��W�D3�Awq0�-��YDxG=���Ub�e�b':���14\��6m<k��!��L���Q��]=��S?]�LjM9���Z�����^�wuy>}	���|���0���*���D3S��p���O�r�ť��7��!>�[fA~E��T0M��Ix��o�x9��)LP&mE�}����-���;S����FEg50�m��&��<���~�tF6�3@A+*�"i��PYS��b���|<Ӕa���*��]��Bfc6��pT]WOa��Xg��MV*2��l� l�Ar�5icHæ����-�1 4a\� m� P�N�+�}�kb�rv/<Y{h��R��.����V;Tޑ]� �!��` j��v��ƶ_��to�����ל�&�ğ���[����O%l������ǭqA������������KBq�R�
%�	@xJ���9<u�i������&�!k�σs`��+��p ��
C�q�߿P�M��X�"����)�����yK�.4���m~G=��
b)�Ϻk�#N�>ި/P�v�6o�$O��u����Y���Dȟ�ʜ6����A�N7�C�5|����\�ڿ��Df!�.}�BNA {�"������HO/	�>�iCo!�	�G�����`�a��%�%6��+��a
�|�NZkz\)�����߀A=WzH���k��b\g~RS���ש�8�PF�ze�.��k<G	���%x>
��y���Q���tۅ�0 cO�~��@����I�Y�0Fy�V)(1��x'0�!���;혅�p�h����*X��:?RyF. �8u��n2K��`~%a#�`���0ҧ`G���ݠ`>������+�Pykѿ:N�s�-V�:xA{v�L=�\�֛��(YoP��CM�_��J$w����ꡐD]�2Ğ���%6�M�ks�^���ZFm��6�:)�t�^�_�>�A]�4��o�9���Q&R��T�m}7e��r"Ҡ���w�즟<kX�b� F5	��Ą5z�EP�Nl�T*�����x���r��L6<� �%	��TR�:��1��T6�
��8�y���ݲ���$��UkB�����Z\z�#�@���U�,��[�d�=c���GB$�!�5l�� Ǔ��#.�@�݁}��VBuN�G����p{ے��b��0�˙����Q��ܮK��*�e��`��Ș����]��#���%�'S�V��Ć�B���{{�\ʼ$5V[B�Bs(aM���)D�L���J�.�,�>���o�%x��8f�T�X%�ʎ삽���L4�CW�"���Yd4�z]t�Z��5����P�#�K�I�_��E�!���cv��\��գ�|Q����L����6P��K�=��4��v[k{4î^!"~C�����ԄN��M�/�u.�� 2�����UN^�_B���.����?~@��Գ����c��F���#E���r4���HC$�W+���&�	\���%Q��/l7f�س�Sey�l�Σ���M7��՛�ǹ�`Wם����XGx�m��UQS�hFOz��L脑�Q�7I��~��E�'tJ�(�}⯵��Y���rg;��)�$2�5����J��	��t����9V�V+�<Q�
*�9�%���1���T�qbqUuGn��j2$�z�����a��-EP��@9p���.#K��a�/�Z@g��JW��'nÎ��c�>CMs��Q5�o���A(y�w�U8���>~��#����9a#�"3����TL��Tq�[�\�KJBa�X�͛Kסp�D���%W΍�:�+V�S���?i���J_H¶M�9p�;���'�0ZOe��w����\q+ʋ�Ff���s)L��z��_����؁��m$�"Cgj�jLW��3@�1i@w
��C��#���$�_�����o�LI�$#F+��(�@T<��K����ލ_]�N����u^���_�4F����=�n�LRaU!�^5��>v�֨�0Hj��99}��{���̉b�S�T<��Ĳխm�/�ԣH�ߪ��ݦy�تi�L	(��4U�(��3�.Y�
 ���
fy�32�&�q�v5��U���!t��)�@}6&�۟��Ƞ8f�r�_�&V��{g"�R�/�L2�"rFkV��E-�<�����R{K��i�vԆ�Q�	��?�;D�������v"Gn]k�S2�|���ZTc1������w,�V��~U�����aq�ԅW~���3=\��Y���2�^,8�ev`�t�����-x$o3���81���Ժ������L���@`�s�G*V!Sc|[��k��CO����9��f�t�3� ��e�0z��p�f��W�g��OKf?��9�	��RA@��*2��@ͻT�SLhP���g�{�4���(��۔ʣ"��ब��x�����c�0��DCTn������B=yE��I��3��s�]�0��zGN�M�J�.��n��B`���M�`g{et���N���P��mj�D�o���#��+���i�h��	*5���	�
�I#r脾����!�X��p�k��S1�ڊ��	����G��3�z'�p�YR�5�g]C��o�q�62[���G�!u��Z2Xи�20-Uw��ҹ���b�B42Q�}��z��R[���|����;�g����'b�޶w;�_G^L7�
�VAs�n��*�7�nAO�v�@'u{e�Xb�g��vm�\���������"�����RӴX��"Rڇ?�?z��æ�鑐]�j7a�'"�9��I��C¹���t��e.@�l@>S����#<-~h�Y�ȡ�[��\��h�:�K>c!$ׇ� ��K/02(�:;�q?Y�6�g���V�Y���'���Z�ϭ&zZ2��oTT@�%�ʶT&w�O�j��ч�zg]�I⡈�k:?������ᤲ
��{�^; ?�K9n�Hj��Z�"G4�]�{�^�_�y��TjG	S5N'�t���pc����uNh��߮x���*B�x�Z���w'rv��ru�b���і���a�z���쾿_��s�.�Сt���V$�6��|&+��(�g.��ª@��Wf���:�v|c[��3�K�SJ��U�=E5��|fv��:��R�pQ�]�u#�=���rm��hs�̶���g�|�bB�?8�$�y�:^5�������߸��YX�>����0��NVYo��t&��L�����眵��
7�@��-��Z�Uuƈ�iZ*+6��ƚ�_$�ބ匀%0544�<�]�MbކN�Pb�$)1m���Su����,��o��" \�d�/�K�-P�)~O,ۡ��6n��6¶[?�Z�g��c�tf�AW����*a�����՞s�1�P%�JJRハk���m�p�&RT_��i�ҝ�0��lq��>�r�V��_�)``ԕp	A��֪`��:�C��r<C5��Kh7VwiV��J!���x��l;�w�P�0�e��V��	�e�b��QB��Q���7W��x"ocS�����J�{�����h���Ջ��$|>���0�~���p��hm��!��L�nO6YRJd\w�uKOy�S��f�n�Y���J1��P�M=�06��`�����¨e��*�:�����?#÷���%J�ħ8i�[��+E�[X��(���yN���*-j�xc��7��E�F��Z�Z���x�����	�]��qw���\� �:J�����֤P��`F_�M�e���x��#�q+� �i��"��.A/'�C����RuĔv�����MFs��p���G@�~WZQF�\=Zg�ߌTv��c���b%�6��i�Q���I�}	�����u$��\��D��^ם��yR��k�ܫ�,;~~����2��S�s�j���&�!��l��v�����˞� ������vl�¼�,����F�ve�4��q��N���|[��>( ��x
֍�Xgm��L^rѯ��R���YTZ�VgqCƛ��ĩ�,�d6�}�@��=\(�а���V�-��#��5uн�1|�Z�e}B����8�v�70�TqR�GD�l�T��iұ��\VHZ�~�E��T��2��� ��'�.�n
���D���~�I����%��0�H_��G��@�f��Q"�T�f7��9�-��/���)�_(W�ln�PdS�rS�}ڸ�WrW>d3aU�9�P����l���y��irࣰ�Y�� 0�XX'�Yn��H�W~5��7E�����Q	9�z,U gZ�n���\����=8��/�zכ=����M8!c]�Т���z��r�� ,=�4���,�`�kh�];�,)87_�Y����^3��u�`q,ꔧ��:������du<GW5��>��6V(�ͼ!��f�*�XM��~EްA��_�*sIrv�QӉ�6�̻��b�F�S`x2���퍟��������l:�1aIZB���{�ώ�:v��k���7QRۦ��(S-��^$�u
�%aZ"�Z��+ÅΧ��ܗ�B�%�e���sg��%r�UJ�i�i��)�si�	rz�
̮�A�
�(~��O���Z!n�ٝ�G��^Z$.�� �~�]���n�u�6�2qe2�̔��{��n�������lF�/ޅ~F�A�I���.K��&5a�x��ݝͤ�*�樏Z��ڶ�D<l�ä�t����� �a<�ޓ3��� �J���4���<j�gQ7�,�u�׮ʜ��������r"�����[wچL�R��E
��
����|���<3��s�'զ%�n�s��]�*ց�#�Dp��D׿��02|q���g4ƨޤs���0�Y*ߏ�D�t��u��~����6����-Y)i����eB=� v)e%`b�}�g�-��;.�;mu>�x&Q�u�X��������� �|��L^L�=8�cX$��(i_HԘ k���W�s�e��Өv������U�GҀ��Y�H�k��6�Lq�"�"�1���Lw�vF���d_�(M������1�����Nna�Ne��M�ۉ_�j�k����e������"���>��30l��r�uX͗�LJ%�udL��'����D���rO�s�'�;��c-*��3}Hn:�D�Sw�g�K�ew�^-DM��t$#���đ��ծu�B�<=]���^xX����M(g�V*�g�Z��"5� ����{�F)��)I��оۚӡFz08�2�3m�u[��(6�Ӿ���7��+xu�āq��Xp�)��2�Q֛Y��c�ݣR/|Y�I#3VA��Q�;S^�/�2�r3}N�%y��فvlo88F�W�@���[���76�]��#jT$���c�^�A�p�/�M��ؠ���7O�*�0$Ʒ��&L���I7P��#a�J��6QT�e���ll�ei��j7�W6C@�����@Jx�X�k?˖	I<8Q?�q�ZM(�-�H�(�c
ۖ�]mts4�-5M�3۝d}�rZe;�)N��3Z��yD��1l�/ZKʪ-������X�1���#�oYQ�W��T_ǰ�]��e�Iqi���ىF����Xp�6���&Cn������6yG�m��9�ox���;	����Y$�H���6�;��h�+;�8��LF�7�k���f�Ɇ]WC=b�1���PRQ�D��sưz���"$5&-i`��I��VL�1�J���\��hV������Y��H�H-g�ެ�w���L��G �r�_���T�e���V�Ц��~���{?�bl�d��)�C��B
���
zk�]IsnOW�w>/\��n��:j�!�b��HKX>�#�R*�x����ݏ9\8�X6~Sj�Yԧ���LzV�ǭ~�-6bFm�I Ǆ�;��#x��@8��"S?m�=D��U�˒G��L�hK�؅}+O~��䩹�ӿ"��.0��FHd��ɄW!3ȥ]�;W6�=�a�t�ᄩrK2蝕�x��J�X)PJ��
)�V��lm0����t�=gLE��2���^؆j(�/��O���J�}���Ofh��V��~ad_�L�-����0���g-�2�C���T�里�I�{7�ċ�1l�Q�{��iˈ=���,�M�a(gR|�������ї�6	�>A�z��2*j��M�����g!.+;"��Qb)��������6j�g�o��ȰȖ�����;��0�$��D9���?���$/�M�6I�|�	f�^^X���+��Rj5�!qOBI������fDfl�tf�R�g{[��d��7n��#���Z���@�@q�c������J%�A���>��Y�5����{�jn�TV��	�g�̙Κ�1#4�"�_����fM�v�i��Al�(H�+Bo̽�J� ��qӻBu����S��]�#YB3`���iͶg�m�$�+�Y`r��U�7�?>4��0��:�8�||�Q���AJE���:�9Sd_k���
�q`>��F�*"����v��H�s�6�F�s��-=�bI��:k�[k^黉X<�`�������6����h>{����3S���i�mz)�I=
�ķ�r�ŷT��`�� ��M2�x�tw�yX��~��~x)fH��ڥ��Ļ������oҐQ�%@g���m��؃�9��2@�,y�}P�?sD��ҮȎ�
Z���y�rv\�,ؿ�W2S��w1}g���.w�9�Z�� �����vrӤ���r��#�����l9�̯���BxǙ)-�ÍڙAuB83	m%��k���q���A��/��l�����d��Tf�4���ް�)����O��++��F��<�a���y�c_�si񡺴>��U�ۇ΅�h���y~�����}N�*���O�g����LR!�H��̚�i�a�|�W��G�~�r̖���#�%�~"�K�l;���^�z'�[��\��Ma��t۫��J�LL÷�K�C��L�9����l���������J��ɣJt~��u-��]���.���/i�p"xY��#�GM�����������PE��~"�,
�%�D�֤g��j�C�^O4�A]5d�� ���2�Gg�̓ș��Q"�o��c����R����?n�� ��KBA�R���e7:�)�bd���W����O4���n�Z#=�i�%�X�fʠ�d�Z՘_, �!O��\4� ӿ%8w�e���j��Eވ�ӂB�*��Ī@�8M\H?D�����7�xV�ܮ�z�]�C��׊�1����}tC�F"xǔ@�Q��aT���2L�p�����F�<�`X��Єl-k�B�k��H`Y�VUm,a��������ȇ��g���D�ZP��*&l1��?�^xic��-ԯ���=&�ʄ����k�+;������*��Q�M�W2u���l.�(�0�a�`�Z�s����P�WD�¬|�)��x��'K�vq�����
U�?��3�!ޫ��m6t}<�S�m��?��_&������y��؂���z���Y0���$��r�!�|�fq�����/~�Fh���p�_-���������ݻ�@H���J���l�[��0�{��)�UQl���y�Ƌ�2�AC��b�.ԛF~>�^;2�v*9�b
P͕i�N��g��%3�������Q+�����`�R(K��W{.��� %�s(��L����Ƥq��]�?�#C��u��sONq�1XM
̣��˔r^�@����Yѻ��@��M$��=;���;m�R�:E;;SuQ$����[���04t�^�b��HVK�Z�D0�<\CprL^�E"�~H���u�֫�wJh݊�,�U�
X���a���a�h}�C�_p����W
*r C�;�̦����&]lm4�C��N��8��!���g�>a�
0+g�bq@�8k�\�"�����AZu	�����A�	�v�(ì�T���9S��D~BBG��I;ln�����-�*�Gd�!� ���>s��{0���̀�C�wp�� Ogȍ{�����c�a�(��L2������Uw�<�D<)�������9��:�U�FtQ�;������H;k1���oҭ��z��Ŷ��:M*�u��/�������,ί�,mQ���(eeg�v��FE4dVr��I��V��8�������d�����5��IG/�d�#���}E(�r��ږ�^�0�<{*��	5�q���(\T$�OQP%]�{�J�Q���	�
C�}9�}`�ǁ;K��'�p��$���m���f���; ���e�<��Խ>��ɲ�����Y�}/�O����X�g�PZy�X!�5��i�dc�,�Zˏz<�'&j8ϙ(�M�Ӻ��x��V�[
��(�	��D�С:-��h�(����7�����K�R�Ց,&w��k*�W8�kX0�U+�?�G��k8�)\w$>J"A"�l>{߯��u5ً��8�݅��C�t�v면Si� /@kf��35Y!gE�ӎS�c��ykw�h�C~Òe5U`r�	f?c ���Pf��� ��=��va�=N�F{ڸ��;?���j]ڊao�R��NМeMr���[��w7�}�Y|Z��Q暽����a� {z�!M�`�9h��m�IvE�6��[�̔.߮��xw�����E@�PQh3;�;<���@L�밁�*��0��r���Eo��Yׯj���6��D��X�h�Z��l���o3ğ����������pf�'���y%���&@�v94��r�O7=u]�n<�����b���Y�]��Sǂ�YF����y�T�|���[W�S�&�_��}���q~}�w?�ճ��cHi�& Tb3��}_4����K����q���p��N����W�b>Yd�K;s��%�b\4n��bZu�mN�;�3�{ˇ?�	r��Ffn:�.��(�)t��5Vt�e�����	�(`��1��Ҥp%q�ן&U#ly�GѲD��CQ�dv��ί?-��o'�^hF��6����_��'�I<mAI��6�<�u�Mp6˃���%��"�<|K���.���w?��+&?�ۯS�\�`u^���T5v��'+��1���u��.+�&[3��E"�hę(BpNԇ��ovl����GO�K�����y�t]�㎗5A:�j*���ʩ12:���8=%䝟]C��G�Y���8�,�mW|����%ˌ��鋸v����kR�����o��1؍\���o�;�����wlI��H��������D�3�*X�����-h�K(�P�u������f��U���%�����gP�$�qJ!�K�����tY����r�ϥC5',FY�^��	]�d3͇L�����먧�˻ɪ�^A��h�#%���"��񖥗N�v��t�#ը?�݈L:�V�'�����R�3<&Z����o��8J]a��A�5�	�էb��������ax���b��G�>TR^����eq^V����6�3V�=SZ�/�XV��+�=�ܐ���]��{M���2��`�R:����έ"�����~:���?�[D�yin�a���mDC��X�`�:O�I��b��M�3!ҷ����I���>w6�Jd�	��i�~����$�<y%�,�G"w�<���!�=V��J��q��GĄ|G�bu2J82<���UQV�19��6k��0�h|��������C O ��q�a7�}�]4$c\��H�X� ���B:��K��J:���H��d��'$����'Kb��5��&6ꋿ��*�0m�L�X�㭊^���u����
�~��{#8tCG!���2s8�Y(�~���8:Kx@�Y?���4��&3MY]͢�RY�pfK:YJ����g�\K���.)@pb�^z�^ڦ_�C%����KI`�V�>�����(�5t6��uR��"��W��i5ƛx�@����AqNk����\C4�� �2�O�2/����ڳ`�2L-���z�픣���gLN&j}-U�h�0�P	Ö?@��;.p���Z �?�3Xe=�4AG�*R��p"���"���3 ��=ΦNU�q�4K�,׷���I��Ɔ�{�u3��JH���xm��H�x��
����a�6'ӽ!Skt,�����q�޵��
y�M����7ٔ(��˵��,Y8�����i7���tIA�����C�qBӄ�K�C���F�D%%��"��(�v
��p@���*)5��4=�h�i�%�!t�����d-���"U��{8Wp�'�-'��Ɗ!dq\;T=D����bvGqo1L?~��h��f�^��-`�oC�"���Ŵ����芔~L�ɶFG���\�Ԡ��'������x,N�B�;�_��]�@U�?���T9g9�	�K�D?b��+<${��\$�0(���\����Q0�0DvL��q[��}��FׯD����K�pg�n��n�0'V���Lxr�1�i���5ƍ����|Ӆ�_G|wz3�v#s��p0T5�<f�`�Lk�$a��|��Y\6�͟�5Tă9Y�:XЄ�q�.b��I�bܛ]�;e$3v�0�y�xJ�L>������:�^��#��u�J���# ����M���Sr��yI��RBˁ��B[&�;����6*!l���1�.k�$Џ!���<V*�$���!�0���� ��z��
.5=6DMH:�	~�y���?e;�K�Ԝ�2b��l�Ff�T�����N��jBH�|�g�t��l5a��g��
�����X#|
��8]�J��������r��]V�ܐJ6:��OaV��l�K�4�uy��(gR�Y���Ʊ�@��ɷ�BM��w����$mрՂ*�s}6�l���UWT�0S'�RVo����|hՔ�!�!���${Z$S����{uh��lտ��g
'5���K�/&c ob���^���(�����
OS�o�w������og�Գ,�q^���#��9��'{J$;��p�3���9Ԥ���ve�Bq�:=jE�E)�B��;bkp�� ������oη�d:�V٘�x`4]�IE���i\\ՖܔN�{,~ْd��k���V��P����h!�kSE����E83�p�,9��PНJ���,{��n�]���Cӡ�nfP�}mǮA�1P�p2W�U��D�B,���B�#3�D�?y��`������K�]J��2�X�i� ���_�aD
�<�'EL��*f�.�ȭ?�Q�����pI�H�1%���j+t���С;8��	2��k���:A�T��:�V��eH��-6w����2LQ�y�jҏ��e�VSry|���Z�W#z&z�i��qz��B�N���/U�V�)��d�"	��̈́�:"��jK4��<��.��)���=�'qdA3iw�|�/��$O�YL�g[��g�Fz��c���F��ERL�`�? N�o-D�aY86[�|�g���҇%TCB��'
#5�9�����e�y��ӖV��1<��޲�����biU9�$ܙ���&\]9�)y�͉���Ώ'e>�Tw'�!��Č��Ϟ_|�٬:��@0���,�tM� ^�#��]�й��F��G�F�C!
LX�<�2ܯ�i� g"��	�¤{,bgI�[�n,ՋU.�1��wH�y�����˲�A�.��c��c��x�`X���7K�)�@9Y˒�����바�N#p[c�����+�R�5�^����1ȑXj��&��-��~�6u<�d_II�.�R�IV�iZ(iO<����!0q?"X#R8L1�Q?������ܓu�w��x��f� n��/�QS,�����k����tOnB��Zd
��aprc�C!e5V���\?��JC��{���pI��C���(%����s_0c4n��gMy]W�5�z�:��"ߞmZ������m�k�Au*u0�~����"��H�������Ь�?m���1���}G���l�_�EF���?F��!�c`�sl��}�A�\Om��$:>���1�����J�j�/�/2�%��j�^����$rk=�I��G�d�vy>����;S��<�� ����qP�>Gs
Ku�Z�KN�	�- �������iWg}�|u�N����va�YT�SLQ��V� ^�%�W��ɗ�iE�z���8E��w��o�J�t]�q+�\�Q'��@m��V�|�I�����}�]3��)����%'��ذ�b8M�I�L�)��]�&$#H����S���P�G�(�өCF,R(��3D��bzҒ|J5N�0�����T�F��1���ʹ5��u�)��N>��ׂ��F�e0t�N�%n��/!:%6�s�	G���r9,{�5C�@�}0���[���h�%�
�e&{V�?�ŤV,���=64lB��[�����th���}	����HӠ>�}��[@�8�����*F�p��e. O�<��e�����i4��0�"�G��Aʀ�szB���T�Q>�~3�0b��ނ��h��"��(��{rsV�-�ۆ��צɔ�)X�J���-�t9PEmo��_�3�AQ���aPm(��L�����L�Mww������f�eS��`c]T;>����)aA��O�MG�C����m�@'l\rX2
�����0u;�K�y�j��?!���p{y3n*�?�.j!1�˅tLg;���(p�O�$^����L�=T��}#�5���\�����n���8�f�0�>��4�bӝ�:'�enO���5SK�IGt�P$�VFB�g�P�m��a����e�B�6ylv�<q���`r.�ј!��E�d��	O)���p�-��=u�-���������}���zdO9��Mϡl���/���1��g���M��yA��g�\	g�B7\���8��M,�����_3��q���~{Ҷ*��
N���Kum+,[�)a�v�$������ث#t_,!�E���0B����
n@w�iӽz'��?��\�t��!Q�6.�(�:<#�agh8�v1��e'$�Tl1� �+�Q�����[A��G�b1��0^�s�V�.�a�k���cYm}.&�M�z����i�B��r/?,6�QvQvB������N	}#���?��7�Gm������r-�E�#�[@}�7^R�:h�c^�	�Z� �~f�&h/�[�<��"M����aZd�u|��w]l�M>�W]&8��A�,Gn��Y���!��BX'�m�6���Awx����m�t�G�e4�^���뇆�S>,VØE���Dh2� S()��,�	�^��yV<k}��� |��y\��+�S��:}޺����
)�y��F%т��9�#�O0��_u C���u0�J2uo����՘�+0��,��1�͟�,�	~�l�
�c����;=M^���� M��P ��F��K�F�Ճ��~��Uu�PCF����oQk9��6�[ՍU�W*Ǉ�=�1�J�����P?+��\C�X,k?�P��6}���1a?j E�i!a�TQWR���՜��M$d�nLXI@�s�#g�v#ە�!&N�
��L8�z�����]�Uj�X�u���5.�����8�#ԏ����$S%�]O�K�B�^S�4�}���Ur�ښl�E�i�~"ل�gS��b�>����X{�����T�L~D/zo��3�b��>�sg� _�<�{-�`'�i�d<�M��Bd�控ci㱠���<�^9C*���S�Z:h�HR����G�[�m�{��%�E�]?�^��<��ZM���8ڼ��xa�E��6cw�Y�p�l_˓4�c=S��4%V�}�dLO�m��n�GJ��8/�|�he�*���G��4���eQ.o������(iG"�d�s?��͞u��`U�����M�Nl$P�
�L(Ç�}~�ȼf����8A�%9��� �����웂��DsżKv���g~���ԩ��߃}����o�tj���\*�e�3����=��V�f��i�Bd�G�a`��P�z4X�����}Q[�P��*�5t�v�?�%���S&U`�bG(!!	�A�۸����+��$/��p�|j���V����w�=űt�H�$E	jIp�L^��>؏0~MM]�d�v���D?�1��꺥p�'xM�����զ�����F};����_)����=f`�a�{K��b�K
�2<�瑪T�${�3�����)Mڤ-R� @�y��hv0�$
CN�e53D"GM�N�M�-/>�/E���PG<Zΐ�ks֎o���P�=؅�ge_��h�u>|�\�jV��X>��%��w����F�ӛ����[�~�������:�I�J��6F�| ��y��4/M+/�*�^&�����!i��*�a��\�{[�}�`�����+vW[}�ȹ����N��*�k�O�Tz|�ip�e�h3�c���^O�b P9�v3l._�!���&�P+�V�Ƀ!s�K[2|!*�Օ.�t8~�K�^d"� �o�ְ�K=�'f��]U}QP�� ����V�o�\�'�y���,	R�h�X��9��U��Ko4�S�~�I~��	N�,�	`I��߈c�1�oon�pc��p��^^*as�r��Z�/|m���>����]:jO����^�ö�\�X��~�r��A����_�����(Hc<'6�~n��~�����e�g\�]L�y��zx�Ǹ_x�`ފ���!�qk:�i�E��V��ѳ��N�k?�T�xW�п�"�P�6֡ �njY�`�ӣ]!u�tO�QC�3��eF�q!�/��=,g�T�8X�Y(����x��bR�����o�+x�`b��?I�pD=u�<�u ���.SE�������qp�`*�˹��k���u��w��{D� c���7d���?o�1Q�o�����FT�]�����F7�0��9�vu���lF�V#��%�,�EwS ����$y�OzH�s��U@�[�3M�m�ѫvqv�!�?'^�AV�Z�Pj�Y��ea�>�"꬏��tt�A=��� 0�
i2��"�yv��'LV�' �T�V�ZY��I��էYτ:>�6�(W#>�����&ۺku��w�<L�}u�Y�Y��I.�	<ۘ����Cץ8l?�nr��dL��J��\&W����6:0z8�%�Aa�����8讑t���S� ��Pt^�Qq `̛��+:E�&Zn��������s ص���1�Y��K�@�vYB�%�ȾQD��17�	�7�GE��v= ���eo'�m��{�y�wy"����Z"�V88	���Drf�3�OΗ=�\]���ʫi�x�]N��ۯEXl��wE
A�˞$��Q��o��~f���>�~��R���Z��GM�$�UxPx��\qVZ�U<�
2����Q��ܪ�'B�%O����l���S��O��v�y��U��v�ڥP��A���uDU��r�{��E�`o=�;̈́v�%D�&��s��jT8:��֪ך[6Uk��uBPQ���٤
8:Z���=��ɍ��6�u��F�u1�=}�A�Ɨ���*��w`��
�<Ȩ&�.��B~�
�%��<����!hw��{�����YJ����\��,=YQM�k;R�6��V���U�K�������Q�Ĥ�Q`��W�9�2��2�/��&x\�޽	��0�8�z.T�Z����Q�!�'��'3�b��&��מd?��Q�c�]_�M��_�>m�Nd�	�@0��"�+r�*/�.�������ov���U�4Ϟ�̣����M~�p��0T�b�%�*B9����8���^X��"�T-jΦ���)������{��� a�%V�F2(�CY�2��x=sM�"�8Tbz(In�:b�uF�[����q�Їr�6��u�9EL�������;�؈�M7mߔY�t�J�f�uo��)gKK��TC�@�p���㗧�g��+�n��I���5�'zN��X�Q��6�"A5�G��ރ�kL��Ė������p_��(b�:���l����(�&^�x%�s�hIW�@a���+6;�6v�%W�HFȮ�,Cԫa;x*�H��؊Ϧ����uqH>v�f�=DY5Q2�q>��{���z:�b����EAtH��49ځh�_f�]�E����f�,3�g�߂���J��-��M��7��o4���g ����=*-�R�Q�D�K�q6_}��t�%�3
�,��(		>�~i`)O��҉�����7���ۨ'��s�*y����+"믰-��Q�[n�Vە,C#�ƇIo/����<Y��>P7��>w�	���4*']E#^`��3���I&����c3l[i�$`����k|��C  �>�f�H�b�/�ѹ��3�
#��`4�_v�v�d�h�x��Z0	&�'�3;�%�����@M��y s;[�FI���tX�8`��̟��b]��d���QNG@sޢ����
a���H1���E�`v~�-�)�\���J�)-\�^������;��#G�0��ػ���t��9Z/;6U�ƕ��yP��r�yF�6��\wQ�qOZ5�i�qv���O�ZC���W�>ls��c�f�=���'d2�}�QU�{���y6r]��u��@�����s��7���,�B2i�V��ߖ;�K���	����f+���ޱ/��d�c\=o�'<�=ɱY�4��h~>�s�-�	3N��M��Q��e�r�El���W�/xHT5ړ�q���|f>�'�窹�S�t��·˶��#`�a�(X?���	���	�ʱ�s�vm%�k�t�\3�|ޫ�WQ��.�e�p���?��~a�dc��9�݂=(	���n�v�2��-����f������.��º�E����:��XN��O�<��(�b4!!�kO"V��8������pŬ��m�]�+ c<��߃�T*1Q��b�qZ�z�NÃ�?�"rm���u�A�:s���H�;�1aɃ�nu��C��j��{hA�xJQU�\#���Ab�?@�u�߲��/#�v@S���]�	^; N���.0�#��2(`9	�\ٲcs6�To?o�b-�6;�b��J�đ�f�lݾ�e�46����;�JS�XH$Q�iR�J|V��Vi�+�/�dR�����a��h1"H�e���+����U����n6v�7;sR~����jZ���!�K� n��:>�����N&��|�jb��[A�m�J	�՛@�RB��?�d� Dwq#i�강=:!����S[\��ʇa+�y93����_gB��︭�4-����s}�p]���\3D�Pr�L��I,�ȯzGF���ZN�Ee��A����à\TQ��S�y<�IJMAHB���0�j��Y��@��,r�	�c�����cΤ�3j \�QR�G�^��)�ƻُY(v8�����<xrG�B�]�>�E��S��k�d�o�Z����2|b�	���	r�|(崚��'����B�o���Ԗ5xt��]M]��e����m{�G��i\o��ʙ`b20�p�5!��o�b�K�5Rś U��qJ���q�%
���kaԀf��RMu�6Fѯ���4�`���cy�9%��U��֤o/q��tzC�ͻ|F���x?T)h�Fz�%ѝ7�:��j��Ȃ����lq��l�5�E�Di��H^9��.,�@�N�m+�}V��1���Ҏ��LQ ��
'g2Un���V���v#��η�#��s�����g��`�g�փ��/����d�p����[C}����H����Ӹ�n�_6�[c���l����s'%ad�e��Z�2�(�0�9�3�	�9I��_ڋb�k�	{t��O>P�x�-cL�<t����y�܈ܚ��v��l�',]�P�n�2�l����,�F�(��b�x@���
I�vh3i��?=ז!:�q�rcK
���x>����a��2��N�lA��	�]L�P&�s1�-/#t�sZD��@��A�Y��)#~U pM�\��4�T��%����Bs��������\�������[�u�����y��fi�f	�v����q�>��ӡk��4�BND�<Iw�U9,m�K%��i�{�_�D�i^~X �X�s}Sǀ#<+^�B}���G�:O�`�;ѵhT+A���N�
�sڀPְ,���o��l��`����.��{_Я(qs��ك��r C��ȓ��)�]f�i������<�PBꊻ+�*�~c�F��"I]|�+��*!o=��mF9��Ի�2�cSO�V�l:��318���͐n�$yf���`
���3��_M���NZ@���c�w{�w�<�u�J0�О](��1���
�&3/���U���,ƜN���o�sq��A�ׄ�$�F��7�+�l?Ї��_Љ�S��`���<oy��?u~òB�v�W��,�띤hoV��Ν��q}y�Q�4�`A�4)��p��?�S�Pã퍑�8N�2B����b���:~�8y��ӻ7iV��E���E~zH1��LZч2�J�_���W����ɼΧ�;�p�WR��Q��k��n�ó�D+�1�&,���������7�"�{?-v<c+Y�1־�}W��)�
���u���Y:c���y������W���C F��t�쭂/�
�Tib��'�zw�qF�� ��b�)1��w�7!X�N��S�n���4������Ei�:���A�$�z1����Zԭ�W��C�����?�`FE뫲M��� ����<��Xo�qf+�ƕ|zZ���]^3v�	�_�G=�EEx�ntd�1��J�"�r;P+Z��И-�B��7������'�R��өg���!���C��hz!.36�2�OAB�]�g~m����	n���o��%<�]<B���e�qJ\bo7�V�0��3pϳ�Āf^ôu���M	CO��t�sZ����Uo�d>8�;&�����E��2�h�UJ��ڍ�_��!�u�&3�J2A%píU�b�����#�ABc�l�S^BFad������G�����,�9�-ͬ�Ch�a�.숊��]�32��������h��)��?4��(I�N��2vX/�ᔿB�����T�@艾3g$]�-���-smt .�J'vGq^���L�x���/�U�L�[n!\�x������ ��!}����w�I�s�f/sfG���T�!�g��Ĉx��w���
f���t����>����\��K|�~@r�G �,�ْ=fg;�yA��v�Ԣ���d����?v0򣾙z�Ha81qx�8��ј�A�f��I��HIa�M�˃�ueF�3gP��vT
l���W�O$墥+�^�n�T�j�O'��5���C�}%O���G9Kd�@�e*sHZ#��r�
	�g��n���a���Ԟf[�ƹ�!��K���l���a��ّ=���ej�.1҆(�8��ܣ\zF�R�m�ءt�N�5y��si�H�	�#koi����\-��{(`�;B�b�ӗ=��]{��]^�/�8 Ӆ���O�c�S鹆��ZV!�}@�2,զjȉ�0D�b�+v�G69gZ�$�����~f��~p�gl����A����@�!)�@�ٸ�r�t:��J�T���
}�����|�&��>�} u�G4��N��A?�2R�����//7�>�9_F V�rzw ����c7d�p6s<����~����N��W�[��s�5�\�����8:5x����T]*$w�Qk�	{0T�����\ K�W���s�0��<��F�G��BW��'q��rV�]cj��<���ұ�����%Z��x{.��$� �br�D�V3L
\Y}�^��ׅsBP��(h�x���Q�\.�4��G��P_!텿�7[S�t�eL!���1	�p<���_K�,>Aֳ(g`�i� z�m��T\�km��V��<P��Qei/@�
2�!�5���m �uAb\r�������"��G��C��<R�$Vz��X@K�Ȟ��Aq��'N��Lpɝq���l5�r܂AQ���C;�p�k�$�������u>r$1kRJUs���. 5.[�c{AW9�]@�g�}z�>�N7��'��Q\v�aou�
j�s'>�F;�3�R��O��A�<ߝI��$�Q�#�⎘��$�>@`�,�R������`C�v2N���lN`h� ���r���Տ3?��U��:%ד������2C
M
`�������z�qɽ�,8��LξL0}�1,Wm��@��t(��M�E�J��r��L���J�L\�����/~�����}��ʃP���e�����f�m^,��x�P�
\�
�y�G�Й��Ed�@]��}���	T�����n��l������Ð[ޝE�y	|���/XR���B#/fJ���[��^P��5 �O�FYQ�G� S�S�k�`CjGHtfY']v��iſ}��ؠ��{����F��;���4vdB��S�WØ��0�/������ǥ�Om.���A�E]F�?v������˶_��Mg8"�|;`��c��~�S�Irt��%T�~�mt��`Z�3���}ί"��)1�V�+77-��7W4p����g��>�~��� �'2�k��K�ʛ��M��������5�^��^\��-��˫G���INp�c�)�Z^���:�nhË������s��[�cz	nt�n���~}>X��75J#�&gwT���������h�r�j:. g�B��݊�sdl���\�GcC�Y�H�i�]��p��a)�)�\��E2h4���I
� ZҬ��M�$ �W�`O@]`�wn.�@ౙh=�����a	��9�0"�O��[Rw3xvs������	�adb���3�}V)B��'i�p�v��F
���&Y�D������Y��$�MP�^��ގ��zpo�j$ڥB����&��#��D�6b������RrI�sV>1��Y6�R���(*�+��~1c6�ٸ$]�Y�3��mf�O/*����n�LV���T���`���0[xx?|J>w�����%���-	�P�.&I������&ͨ�P�l�0EBW��~;���*�����F?��L�}01Vowؑ��c�3h�#@�q��dO�v��d~~��o��'e�-���><���~U��֍����>3VZn��V���n�+3�(�Ђ�0�8��=G�,C.7��85��Q��Dڊ���:)���"�m�9���W�F��ޏ��y�Y��E���O�47kOpm��r��@��N��`�@��#өxRT8������qnI��i����_3p�w""�O}�O}���a&r��`���h�� �Yt%�^��Q��9yכ,,����L�f�]�'8<�\ (��U�jQj�m���e˼	y�*W!������M�!i1�L��k��]�^�!l�t)]��ѥ��u e�A�n��7d���8t�r����v�8W�W5/�;DG��L��Ng���(%4�;�ٰ�6���xi��$k��k7�ɕ��~eדQ{�&_�1��7Xh+#��@"���\B�
h���G�i��	��k���S��
=\��j�JɁ;��x�L����|~�̭H<X�i�a����P�5�C�u9�q�UK%�dQz�$}A,�\�*�L�Ȳ�l�H�������ť������AFa��H�ff!���\/WPz�����*�W��Y��Q�^	����r������mR�B��@��\��4�h�#ъ�WK�f�On����o^c�U5��`s��4Ij�xs4GK�t���)�&�/�S��Fs�Eh}֋ҁv䖃��/Hhr,��o���^�Ͱ�=����<)����^��g+M����D��-�,����8�,�����<�2����\�Z�VC�)�,�{���֔t(�����2ȗ��E�����q.a��V]�Tr�֞ΐj٨(��Ϧ�Mi�!�|QnDIghޔ�fl%��/?4����gr�����3�L�T���$9Ù|�gP��Ψ��Z*�+�}5k�`��R�u`�Jk�;Ȕ�1�ס�_��<�	�w��ך�[��*��J8ђ�^�J���(󹫨a����jφG?�$�3�m�M���22�3+��9�=�L��	qJ	M_��JgU߶�º�_�T6T},�X���EJvDqs��(K��m�Q��rtfaR`[����E�%������{wCa�fc���C_�PC�-�N��>�[M�R�v�70C!��.'S)m�����h"TzU�V{-p*&W�����)2��Y
��!j囶vR�r��>�Z/�_U1*bT����_�(��s�X���624=YѼ9nFO��� *Am�#7{���~5ݾ��:]���!����NK��K9�k�"V�=_��e��}NE�k�U�"�CU��-�cY�ſ�J�dY���[p^��y`��� �� 35	��#��_�5�G�\���x;���l�,��/|)�&���:��j%2�AL��ύ����̇q0�/��>5q/�*@��t�����?Ds��&޾��v���ۉ�d感���Qp"m��D�P�"���}��c���6���#��t�+cɹ��$�K༃�O��:ȳ�"4%�bgf�(�����)�F�U�ʘ
.6�56h$.�B
�m���׺����Ծ�i��,�j���ܮS�V��\TߍUFx�]Oj�=��k<	z1-Y%��aqa�����q��������$�\����dr��0dQh��W��]uQ��B���__٭"k܎�]�}��y~�.c����'�^ۅnN�sح��m���F����O�_�y�d�����]�
�"nN{ʸ�y�&~����OY���	_�����:�w�"��QjN��,�x6|L� 2��٠���7
�R4���+�#��?{�G@�ax�hi�fqWK�u�
%�
���J�=�{g�:&��́;�w�e|7:���K�kmz{!�4z�N���0S���
7le! 5��T%�	X�TTl�Bs_p�@��ZVV V!oA��O�N2�*:�"�X��ĖM�$)�bc:�wl-��Ѧ�W���?7|�)��]c���� � ��А��|�wX�j��~���pZ1y>�N��8�r]{�����,b`⏎��=�/�\ީC�mG�E�e�M-��B�c$ou�<�����K��⩰�d�]�Z��Hb�I�T(����2�=]辄崶�'����"Y^b�s�n0#HG�J� ��S|���L�pX�i�X�
�1� /B��Ü��J
G|�^~4o�8�?�݂��|��r�C����@��+%(n�A� $��^��Z������ۺ�Z��D��<����EB1�`Do�M�=oB�v���	���?5}$�PL�P�w���~�	�Tʣ$�S��7�4��-<c��t='�p��{�I�����%��4�q�/|���G=�)����z� �GX�u�9ym	) ޷�Cn�~+q$]���{c��׷Ö,���G��ii"h|��eG��F�̇��$Tj��g^��v4b�H=+�ޒ��͑��e����@�Q�!��L�o�,������*/�Z�J{����?|(h���ԯ��!���G��d�q'���z38��~�`�Zւ{H�����ו8�E
�a��<�_�%i�v���sn�����H�@u�y파�.�s|A�ݓC�����'�T�,'�CZ�]�-���#7����a�U�b;�7�o�(j��j����%�aP�,�x����2�8"����;�.t����NO�=�/� �̄X��pԏ�;ZB��K1�D	�KԐ�/y_�@�<���1~J�؈��x�C�Y-^Ȯ�J�<���s;��Tyzy�6�M>ۥ� �!��2�FP�Ϭa�ݭ�Cpgg�w<zh`�5M+! D8.�Ds9��-�7��\�&3�ǉþi�^�m�b�_nHL���4Z�`�	6�E&b{���I>�ܑ�O�F?4>�ו��jk��<r[�z\z>�_|�?�\�Y�o�����5��3眒����O���Ȟ�Z����}E��
�0��6R�[g6�޸the�)�2�\�f;�0�e\�7,�@���1���VNT�U���drn�l�Fv�����OB�jYd0��l��b%�UX �3m6~��{��
J�D*���.	bbB0�$�7T!�w���F�(8S"̝0�i�L5X��t��_��΍}��X]5�Ч��͹1�E{ ��^��lt��`�6�@14�8�|���8uvt���?���f��]���	#T�����, r���O��D{|O w9��F_&Hm憰K�����b�w���������M�sW�1"C��>�
��C��ko�P�1k��	��4B�!�����XEz� �b��@1�d�am���d�!��^�E"J����2#��@׏N��[���T���	��9��9��P��BZ�t��3���{j�mB,� ��	@S/JR���֘�^���Ť�������!͹�&���7+�Uf�?�5��!'۳c~���S.���*��aV?G��1��Rxa�zVM!����l�L�I��'Ub�6�\,����S�z�9�b����K+����(
8�RO�f#��b�p�{�i;�ܖ�Qt7K%<V6܆,y��E$�$`���r�Tmd��<�����5vh?�wM�&�(��^�&�����z�m�[���L����%K���L;@`�[r��\�5O.�JFp�MBF�B�y!�,�g3|�O���-|z���e�c���"��2C� /[韉;�*�f�uO��E�Q�]�@T�R���l�$�ht_��̸�M���AG��Ǳ����G�p�%��o�<p��߷ E��E[y��,Q<�VZ�9KRɇ	��'GoN�O�M�ո�:4)g�l�E�c��Le*�2�a�����z�_IE�����K�씈i2�&8��nG3���>
��؋�- QV�4��Sz��!��aq3�?��+٬�Tǹq�o��ɵ.0���M�b2�aX������巀�����j��n�/��psg����Vslk�2�K�N
؛��z��=��6%�Z,ǔ ���c�����s��%�`�՟��M!�
�+ T�5�z峉ftզ��ݬB�;.���:ӂ���W56�e�X�%��!�����;��mO->O%�VL$���R;��(��^����K��N�|E��Ck� ��Rq����ڼo�*@kyʿ�S�E���_V��}�����jT	C/;G�,����S]@�����/<��;�~x��}Oom:�gߟQc!��G��� !=x��M��Zُ3gfem�L� ��|�c�ӳg�a���8�3�T�a��&��f�$8�eumE�м9�������͞���l�8 ���'۾��#ٖ�?����అ��E�#HT�zA��.O7Pp%)px$7(�3�%C�VA?Jsw�+󧋾��@� gE��<��kx�c�w��b�>�8<�o�
y���F�~��5"�-?�N�p�W�V���bq(E(4���j��y@֙�6��Y(���^=�)ꍵ��G]Q��Dc%=��f�� ¨�爵��s��m��(��^A���Y��SCJ;n��ݍy-*����#���3�6Q%��~�ӞO!�\��Vҵ�1�m�<�vbU����V{��/�����%ܮe~�����Q{
`!���j)���ɫ�qU`�L��`��v�8ìm�Ig�n��2�L����▗�<V$d��z�]^�m�Ug��l�'�J]�����ػ���9��Gζ���4��8�@��)���ꔚ��)^ݐ�)ɇ�\��y�F�[�`3"�I�k��h���C-&t��=5�U4-uq	1�،:~Dq����bS҆��=$i-�S�V86�WC���	����j���ݒ�~S��@�l��Ap��vZ�����������TH�S���������~a�	�z���V��_�o�B�����-l�&�
���e��?�/��a9�S�UBc��ۜ�X0yf0�׼�����6�_����#3F��;1"�y��IAf���
��2ߘ!jj�Z�72��wg�,����"#�i���*qcY��hi���./jN��!9�e��n�e��J�ڜ���8���s��<\�i�k���V�h-��c���f&��A���k�gm�~�:�$��D`2W�.&�'}~v��#�$k�U��&H�5��ÿ$Ɩ�H�����O-9�4���n�_2PQ�{�v$]� �r��
2%�C��!m�Y�R���I2��֫|ҩNU�pq�~:z=�b��?_�
[��ha�.�F�ߺ��r-zE��?�����9�=�uE�_~(�ŧI77K����T��^�0~}l�$��w�����ހ�������Fة�U���3�I`��vH�lԾ�y�rs���@���(f089&'|�O�?�߻ ���BY���jS2ѓO[���)��(��J�A��\���
Ӎ����V]@0Sh@�g�3	5y�	�u}��ʳv���H��Hh�h�<�Aąv
�߱��G�#&/��5Ӱr�f����t��{.�zѷhh
w�಍�H3cx��1=�Y1����ftE�%B����k3R]�ӳ$��R�H�	�N��NW�:9��B��%�V�I�+����ZTғm�Y����.'ut�x8�v�r>^\��h�0�0.V��x�������S�T�r6��.���paE��9��3�~��D��܃P>�n$�r��:8I��.�OX���I��T�(z��_��}�A��~��m_DƵ��\'��߳p=`{Y�U·���2ˬC5c�胢X��!���(@M #��O"q����@�:>������о/aa�w���G��4��W���-5̠���`��0S���Q��b��Ǝ���}�*Mߌ�`�܇9Y��"�D3��N��J��J��8�Q���BzCr�	"l�	��H�5l%�K�3)#hA�ޱ�x�L"�r��wcO~3y#����ׯ��� >�/ؓe��+?λ3��W#u�Mk���u8�O#��5�t�
���.�S?�Q ���0�/>��|��GrK�����T]f�3����#f����"p��8W��1�=e#s�9F��2C�A�ݩL��컴gy*�̔A}�I�. U�Zr���*1T�|��9�P�4��cW@�O{l��kZ�ϳ�CN��wyhJu�*_k*����e�����	Q;���].vHC�H^��� Bb1�Ĉ��|I�����@c����$�^A-��XaV*æ3!�li�{q������U���g�1≗�s!�N!R�"Ga�j��G^��[S����M�5�~R�� c��|����
��y2.�P�S#��ǭ)p1H��m���c���Z�bA��q��d������t�2�-�(�5Y�hHga	>�����#p����y9\�WcOY�P#���אIY~�G]Q�A���q(hz��?տ4L�Mjѩ���"�e_*��W�Z�I�{�� ����KbL�cb� wa��uo��8���21���gBr�	��\����׿!�}�)��3�QR�W*�b��ULwWm���+�i�2��]�=E��ű�$�s�6D�OTX��؆�r��>]���m2Ќy*S�&*+&��*R�_Ff�_�Y���Ȣگd����Z'��%��4��+�������AOC�2�{�.f�~��_�\-�)�9�5 ��w�eO���t������/o�ϻݾh�>���
�<>E%�;�n��uSx9��ُ���ɤ�=>��?e��5��_C�VN�?;��Wt�^S!po�u����u��K�H�5^0Ⱥ�A�Q�=���x�a!��f�|���Z�����t�nߢ��$��b�3�oO2d)�*���-dMj˵��9_�fz��QT}�ƞۇ����gʞ� ߒ/G1bV�����^���ōY�;��ĠĆ�Š��xe��2��&E_"���]͟� N[�V?��ay����z�����J��8������&�#�=kwD����5Å��_F����y�5?W��E��&ǅl�X�Cȃ�p���k�a6P���o��[����K�Q�MU������K�R��,]3�F�����<3Uy)<+�l�4��sJ��VjPvS_��'\�Fc�L,.��q�������a��g��Gef���L��"W)�[�9���/�lx3�����"��.*+AL/�?��n�~3e7�~�`<���
�����\ӻW��(o��m"@@ő�MⲕxW�˒/��G�Y��h�\����V�3�S ��4�Єz�H��ۮ������@'�f�@[	G���Ւk�q�!�h{�ک��#WF��LףWOF,^'`�t�e���ޙaX�!nFɈ%�uܼ�)ב�����0��h9w�+p�p]��C�D�����I�Ԡ���z�j� (�mWHSEP���)zJGׄ�Y����W|�j������8�Ȁ�J��n"���W�U��Z��)T97�sG]1P��~��1ks�@6̷0SU�t�7#�v3Ǔ�ϻe��j����2��%��6FĆ��.[k�u���O��,�c����~��˾�IfK %i�s�� ����E9���R	�kј����J�:Ei!���[�~΀��ga�M]*��H�ޣ|�t��Z��
8����OGAj���w㉗~���f�5�Lk�!	'�������1�f�Z��h(9�Ԋ&�+k�b���W�ĕD���V�D�|!���Ɍ<%֫]�R�:�>]A=�):߬��x��|�2��PL�]��W��<KB���<�5`'^�J����8B}i�ka��ٸ�X1',�sN4���&&��2����p
eW7)v�X��uD�Uߪ ]�=#�������[b�]w������ �@�1�f�<0��vJN��NE^;c �ٛ�L�/ ��;%L����m�f��F��t�+�`0s��wߌ��g=��`�S�8���*Wݻ���l&�� �y���+�]����E�c$����>��fj��9-Ά��:籄��Q����U�biq3U�M|�T\��R�WɁ��`�F�|� ^��^�L�|�$���QDlz��,�Ѻc+-�N�ҋض�8��8��3����#���B�W�P;|#�?�u�#�O�47k�y�W0^'P���EuH=<�S�,�LKf�%S������ƌZC	:_PIַ�� 5ru�nI=U��&�n�=(�j�[�u�F�Dd�t~��J�� ?�P.��W
�c������!���[�[`3�׫|xQ���=�&=B�z)Qj�hO�m�vj{�U�b�q$2a�"��XK�dp�m�'[����np��c��Z�-R�*`��JQ�4?M�-�nA4��<
�Tm��_�^�� olgGu.o)�c�hv��?"�6�T��ml���w�4�f#f����uu�3��1�T��o�T�N��F�@�`v���{
,��2�LY�TՐ9B�lĮ���X����C��������"x�K0����a7�
���r����������$�N##d���3[i�/*j,��ǔ�������^2�"��^+i����Q��q-����>ƿ�發���2_�dRf�/�Ӫ�</#�yK���Y��/���]4�Yѭ�9��i��S��P��Qr���1�:O��_��ʗV#%ʭ��ǘ��T�K�)��Q�.yv��H��wR��4k���Z�K6x.պ��i����u�Θc�,������<��f�5���D��3����=��5O����O�n�HP��r�0<�|JZ�ZH�� 3��6g�M�淮��HQ�`��a���j����J�K�t��5�6�6+6�{�/��o�*^�>�#*��w �Օ�⪙�Z�P=��_q����H�X�Lg�0�p�șn�ls]�o*��"U-���y�O�@����Ý�2rB%���v�q,��@
�Ǉ�("��(>o X�2����K�>j	��v�WzE�|"
=f,/�k���D�bv�3���V�l'cN���dG�ѵ�S*ȯH�ꑽH��d�n��:���Q�Cas��߁'��G�W���_r���|N���#�cd�쀤o�L��W�2����j�ygQ��z�.����k6i������o�ʞDa[�V�*�@����:(Ku�4Kh��(�NjV�n�s�#<�Ek�K��W�fx�����Q��)6�6z�j�S��L_S�����q���]uf
�����C����`A�"��[nVu%@�t,���Ձ~�S�k��A��.���nf���<��{�74��M �6"��Ve^ꢄK�jI���!���c��zo��>l�����

/ܠ	��-WF��(���y�����%���#>
�?7��Z����K��}\�qdL;�R���4�����Nt�J��Œc�ݾ�������&u�����m��U�K�K�Z���,�ni
AD�5��rC�Bh����·���yeR� ^�q��Dͪ��(��x���טkg�0��Գ��gpBbr�h͜�:��(�ve`�R��%˗�J;�]��!�etd�YL�nI>?�vuЉz���#G��m-Ď�(�/]����*Y�>V!����@ܯ�j���\�2��U{���>M�s]%�hU-����C`��MiԾ_�	@�j�2}�<�}ⴺx7Z���h�8�'��u��OnP������d�̖�["�fr��ߋ��<gV�i���u����&�"����tdp��~�˧�Q��y-����m�HQ�3k�hA��pX�V5q|#e�(��/tf�o� �7�\�4��@���V��x�p[�}6fE�$\��GUM�_.��/�q(�����*�������:3r��&�1og�C�"�����RhG+u2�?̳,���T鉪�o��	D�N��r�2��jR�K2���xr��|�H�WU�7Hi�}�y�ޤ%��2��J�(��Bث�d�VU:�(���|��)���˰��ؔ�Co
!�[g�'{b@Cx<�g�Wmj�Uڸ�1Ӟ��0f4�_�U����U��I!?�Y$����X���|���6�?;y���̟�ց�O�Tӓ�V[G[�/[��,p H��Z�1+��xa~|}��]$Z�;�l6t �^�9|�O38,d�'�Z�E�'xN����è<��f�+ԭ��v��O�-!���;���p��DWlܵ�8cߺ�$�;� �\�M��N����%G��oX4ݿV�G׋��� �6�+*�Hg��^ *����R��-�y}�g1#��
+}�H�X�\�9^A{?����E����yy���5�����/��e�����5�oewY�I�7��"h��G����*OТ7��r� /��J���(�����o��5+����y��9�~�i7A1g!E�W�DBؐ�mr��!���$F+Zݽ����
���׷Y�O'"~g���� ����g�`|:@(��A�AB70��JM�10L!����� �v��Y�k����|��-���h2i���6����R���_��F��D��4���&L�/"y��1}4��k�ٔ�w
l.��R�|e�r�
�ZM�!C��&�8�{��Q
�i Y8�Za��r,�eG��5�pb	>92��f�^�rE�C���+�r�h���H	U��M�����K;ZH�{�?�@vey2�ϠD.���sr���?��k<������{?�<;�'cH�9w��"� *uǎ���c�  ���Z�h{'�1��C���\�wyM`����;�J) x�9<��:�IL��Ⱦd����ڮwD�:t�C�	g���v�>�(W[�t�W�(eCF��;�eV_���J�uנ�B��>^���n�S0���G�4��t�p�10�(jsg�R.PV�/�]U�l��;$l'v TP�j�c��8�?�,�^c%o�<L!�^������(P��=�P�%�Zc}H�^�~N#s�ė�<@�e�|�Iv�6R�l=�{L֭��J�� ��:>L�o�r;P�ܪ}�vBڢ��3��V�t�^:Z%xy���&�"x��R
w�i�����Jz\lt�u���d��i)�~�t�?�p+�x
U0�SRK��o��N�C�؃�n���!�/3�8�vL�Ad�pU\�o򨩷��'OD]�O3��'��)��s��~�iNam+`N3�hs��YQoԬ2��-P�ҷ��wQw�`��HI�X�Ւ���ĕb6�Q�X����D�H���`��N����qى�T�j݄��D��H��d���j�&��m��������f@ ?��dn�M`��n�f�6h��uS]�;eaYH��l��n	�WU�`��Տ(���^ϔ��I�șx�M���[T�<�_��� %��3� }5��E9��o2�]��c��}��OHS�2��D�4O$l������%�L{6H$�q������<g�${��&��e(P�L�NM$����Z����1kk��hz#]��%��}�z�Q�tFeb��	��)�W�*��T|�'���n�G�cDo��������A����|��j���jDx����r}<�Kr<�����ٯ��^�-��d���+�rme~���"�mئ� ù���|-��Y��������� 5�k	Nzr/h����>��,�̝�UϺ��?�z�Y!}s[����r-�� �ٷ�4���z��|��S�#2�f�p��WMA����>p�M���X�]
�=�n@m���4�����mU7En����3��`vA����R�o�Q���۾a��B{�2��iD��7?���ukM�s}4�	��;&�ϴ某����ϝ�V��f�Ů�Q�u9��߱L5!�[�� ���/!��=	�De�L�����ݲ��3�����l�.u�:Z����i0k�����MA2��;�/(u�e�Wf`P�_��.���f�v5+�??�рJ�0|��e�E}(��(&�Z��O7���bk�dvt�B(R��iP�&��ɟ*1a�m튧��	^�o!��Ν�g�w1�í:fW�7�0�wz���$Ҝ�]j%m%G��Фt�௉I�u��yU�7��G�䛐��L��r�ri�B�º�pW���(���������ȶUa^?�O3��̷T�=Z�����84,�%[|���J�_��B-�4}��O-�]E�ä��_4p��Ad���G���%����[)&�Je��+.����w!�gf���	�X�:���5����jZ��}ȩ��􅼍��Č¤��S����@��5#`��ߟVdj��9����?�&ɮ��"�?��������D"�<�L���ӈ�<p�Zr�t|���'hҪ�#�F����:�J9/���ǥ�s@��@$�ԇ-������x��Yt:��&��37��Tİ��^ ��@��q�עi����7��z�����3J�ˋ)��eR45��a�D���r���Z��`�҇��d�I�͔�U�Ԙz��8M��?QCU�H���+��)j��q�X~@]�n��=��|��˙��.M�eh����6��t-P��z�ϪyZ�$�́�%�;1�d��P9I���R)��Bi"@S�DN&���k�Ť@|j�g#T����<�3��ԛ�6��?�
U���`\G���o]���cyp�[[lfR�$-Ε����Z�L���(7�#��m׳�5�ۋx�}v5^��]z�Zĸf��/��{�� &�p̝�J'��Ɍ�-�e��ݭ��L�����Q��VRn����e�����|�u��c����ղ�!f�`�2v �l�����[��Oc��� ��#�e�Wv몧���I7lϼq�T�d]T ���cR=����[�	�F@@�d'2ֈ���'ò9&iX�k >�r�KQƲ���1mJɶr/�f>$Є���z��.UWz�����.�����⡯�T�/�L;��mb�F�Y��̄��^a�F�rf\�4�Mlt�z�.Ֆv�KTMT��p�
71%$�6W/W�J`&,Z���&��^Q����򦐐W"�l�)�[I�&X�SS�����4��)bl4>m����{��Dl��<�_R��7$���Ή"πw�-�����}�%r�e�ca�>k����|wsqǭ&X�������!f w��+F�%���(�W�Z��+�h���J2�MV�P�:�����7w�k��9�^�xCǜ5�8˩	��<�8 ^��w�=]P�4B�� BP:���2�~�v̍���+B���z,�N��bڟ��#׎��֛�\�%�_)���f?8���`����o�l���V�t7a|�u0+��m��XD=����gK"jy���Ø��n��S���ɕ�+ҋwI�����~AA� �gil�zdۤd�P�D��;19��l�������㵲���0�?"0N��Ym.�"��J���B�k����O�[��ʺ:ةco�z�o$���+� �����\���
A����~rMMgHM>`����;��L��7u�u:e�M��j���� j�����GÍ���Ï�V��[(!�\������s�גy.����)�,Mt�f�"Z �>�v��'�v4_5\��l816�-^�A�5�� O=�E����8���EkD�~��㥄0��An�to��M��m�/��s�<+t�Hjq&ِQ8�F�&�����NS�����#����_�PYda�|����M�X�@'���y�R�WKJ��=�K�UVs�8%��D怨 F�����׆�
�G�������ʀd�6�����A��;"^�&%�N�Q�
E�F���H���Z�7صX�0ތ�C����*2��	M)�皐Sf�m!8=7�SN���'7T��/���-ʁG.r�D��lS+9XY$ŵ�$^�����U�qï'��O�8��^�I���M&���������s���:�K#�>��Gd1�����	�?~m�x`�Ѿ?��yH��ŗfQ0Y5LIٗP������XϨ��$�-¶�H2X��w.z�KkU�ݎA_k���ƹ���	H�q���φy�|��@�J�tᄻ�Ef�ۤ��%r-,K8�H)jU�:u@1�E�K���Tz�w0��}M,,��[�~�}�GW(?\Y�1� �z�]��B���GHz��|,V���Saa������1�n)E[�.4����_�{��x�2��}i�����v������:^g�j��4逢N���5��5X�����\�9�u�Tu.�F��	O'h˝<f���\|x{+�.�m`bˏ=��@��t�"E� �:A*G�S�Bs���y6�?D��^��2Z$2��9�㰊����4�y>&__$*!��17�n߾���7��x?���Y�c^�����Z�nQ��Q⚜��փ?#��$�4+M��7J��+�v�'?$��t�3iB��;�	uZ�1'?۽�a�3��ь���uP��g��D�m�OP����9UiƘ��4 XZ���&���[аb�G�%W=C�D��sh0���!c�Q�"�����H�F?����Cl:�~��X�)P�0�#��O��`z�\V✜�����bvC@|�4�j�T�+������c���8�W�-��3�"#v�ި�wZg�,l�
/�C��7�k����2���`����+�e�
0Z-���i��$ ǆ�C������GwA.��Ew�_0�(a^#|8��3t:���f�N�^p��]��r"tfv�:��6������3��8Q ��r�00���K���8�L��6? v�*��&w�l�]��M,֤kz�u�K	�B�����E�������[i;��q�&&�vs���Y��1�����������T��K�8@�O��>���m��k�E���o�1\��D!�Eޞ@�^�W���ۤ�m�ʎ�9%玲���;<�C>�_����s��o�O���7���
��ћ���O6������uw�|�i�/��g��X�]��۟�:��o�x����x+� /5?;��_<��/Mf�hi���H(Cvܵ�̄�GQ]�HG�:�V�����x �Q����µ�F��E�R����	yMr�W@.&�=��ĩܓ���Ѣf�#q�[gfu�(�vdX�f���)Em�S�6��0t�*d�N�,��lK�*棻c�L�N�AE�'��U~"��E�Rh-~Zu�����7{"V#YNHG�8g6�b�>b�^��M�n���+�����`�&�z�-�����3ocm�)��,�J�U�{*�Bzc�"Ƃ�ok��O�b�7&z�s����+����HM�^�PF�k�.o;��éӰ�ǅ�4��P;�X���w�]H���)|������
}։�'է1i84������I���萉%8�� �tt.wX���#���$�b$V�� ���;�����Vb��ʣl��Gח�!�`!�I�K�'ߤ���X��.�:�>�:�x�/7¨�%2vz�/I�G��h���]p8>%�Ĳ�	~�ŉL崾�k��o�u%a�K���dA>��i�'���&����Nս��ki=Y�E�v��h��9��)�.)��]'H�Q��/�T�&B=�U��d�C���������w�Ĭt��bpjZ�m�`��1��LF��m�,8�P���޾�)���M�T,KB�&i�֫b�@��	��5NW��L{�zQ@n #̌*��;�)�ʺ�C�$:�4ƒH{��ɹE��!��i�� ��%��&\�%�| ��=��1�iC����}=g�0�ɳ&]ӡ�S�k���2{`��À`����V rL�s0�+Z`�̹i�o(���}' ��3���$_w��zP<�����>UMlg��H�]�:�j����Ñlp#�Ρ��&�E6{q�/���w�4�ӏ�>�xM;8��Q�j�����o�9˔<r�'O�Q��)���Q9��ħ����қ��<Z�2{53Z�ˑ)�ö(|�;�T�'���^e���x��J.�D�z��b���,�����5��B��M9XO˫^���'�j��㊇�>���/�>�(|"�s%�&�=+�߀6ŋ5&����(�p}wb�ƈ�@8��[�a1|�:�;�=v͜@�24*\����ء_�ae�a��Cl�⳦N��d͜�|gj�͹�<�E+�	TqC���O,.��n�DD�������(R�(�{i�47�
����d�Zj��^9Wz���B�y5�K�R3��/^�#� �/�A�,~.�ֹ���J���ծ�H��Gv�V�3�rr�g�#��W����F���L�9!��\�E֎��"PR{���7����_-�h����ad6��15�]R��FoT�?���P�W���3G���Ƅ�}�CW[f6Ǐ4��
�6��A�q��Q�h��3Y�+)_�!�q
LT��RZB3����{eRd��0-�0��<���m�Ϥim]�y�Z.;}������9<>��,5
���.A��zptѻB�؎�6�c����Ua���:�"���^E��@ոR�6����x!�͟�Ghh{�r�~Oo�X8�F��&��yz�6��[�1ar�$Yu2���%�c+mS�:���x��s��A��;Ԑ�g�%ggz�p��I���:O��D�S�s Y���
[M�wtb�N
(��n�'w��
��d���z��8�\ʄ>\�4���7�� =Q��Ā`�F�F1��/�
�)�<#�8`j�G�E��@?��oC�_����&��"���AI�/����wįm�}4�j��j�lo��W=m3�
͈(w$^�ƝZ5�c0s�~ĭ���Ak���)#�Y{z�0=$a:P%�}Q���{�o�L!zv��S�\��ȈM�ݵ�8*{�|}*hp�wG�q�Ӏ�ݎ���TD�N���2�ᦧڧI�~�fNyl����␓�����ø���56%�}q�Zs���ɠ1[�mx�%�_(b�����bi�|�>��z�T�}���}o�I��*%Y��	Dp�N�e�B�ː�LP�)"������|���U^9|2=S�����m��*	��S��iTKMQT�L�gp��'�ޑ���m�Kg�:XM�.HYg�3���O��CJ="�����	&���>�x�3���˩���&�757z�;óP�@���0\��~|Y!������;�	�cv�K�i������� ڹ�+i!�����-��fW�����"�n�+�
먙�i�[]��eH����fE.��Ix��B4���n�/�:�_�Z�"UL��gK���xl�b'v�$�C�M���f���/�_��@7�y'�2�*4÷�*�d��wb(2嘨��E�3�+1/㘂�y����.vWt�R6��NӲ�O�dOD=�(;�����K��ja2Ug��v����R��=<-M %�S�=�2́ݱ��� �DW$P�M~�IFNm��^e�����tԋ}n7�{�C�1x��9\&��U�լ���������-�cD����7�_��CE���¿��	�;>H�@,a�=G�����<@���R��6X��0j����!��1�=)d�K���9c��?{����o���f�jژK8����Ô 2�U��YQ%ݶ_Pv#�h��j����N�
�o�@v��8:"�W������ЪN4�\ {h��v��!h#L�"�{�{�@h9��r�vu�MM��ml�+�Nr3>��#� �K��:������&�/m�i�]��`;��W�3���n�y�S4=́��c��+�A��I���T<Hy{�^9�B;�ɶn����S�e���յّA��:����N2z�ԥ�^�)����8e��B4p�!⚀��K����X�q�Gjw���i�w8c�^��Die�����Y.>ߡ�x�;�l�OȐ/�MR�`�M�����������Ëh�9��Z���;���9_24t�t���YP�=#dT%<7��<Շ"��Q��E� /�>]���Gv�t���1	�;��&�)�tA��
By�4�K���w��ɌR��F�e��:Ҧ$c��Y(Z�H���P��?�/�؋wL!��*�UM$ݨSu���"�P��$PD�k���D�&�)\=U�u��Q��x;)��r����Nh�w5��/�^k{�¼'��6�AA��J��C�z��1c�gܖQ'�|_=��o�NQ�C����X}6w�}3��u�r��am�@[;���	�n�⾛�\���N��9 
I���������[k�#�D�����7ፕ�D�0Pj�m{*ݫ���(�U�x�GC��F����f^u�Dʵ�i�P�� 	<�&�N��b�
�,��7���;�,�eRWN;���@ˑ71�I��(7k��1̪�-)3,h�yI�w������O��b͆Q��!����=RKtx��$��nP�X0(��\l$�Xs�o��8M.���O����ඔ���4��c�Û�e(�E��2ONό�����l���ە����it܉ D���I20��HH`a�&R�ذ��K+���m��H���Z?�>�p��.�����C&aY-zP���ʬgfӴJ�K �l�Q��ڶGU��s��~,v`��� �Vc��E�C�19 �pREӛa,$"+�Ŵ�_�yNT��1YE̺A="!n*ε�� �v�>z:p�cK���A��f�ԓ������+���ߗ�h���;ؘQt��BB&{.c7��l���`ڃ� �_��C5)�jF�1dP&���K�������1_[�����:;����Aia�NaEƘ�������p%�M
�ԊY�U��Ёɏ�J���j{8}#��������c�,xa�Ql�`�b�RF�b�؋/3���u��{-�QK�t�S�.v_��.tf-�g�E���$�<����N��%\���d��a΋_Ȥl�mH�+-<��~��Ii�>;�7l)�8"�:kZ��u��9ri/Q�6����S�F oL���[~�1�{���h�����{ҿ8�.��� Re1��<�>q&���خ?O�+n w)�Ŕ.㯲�\���n��[�e�.�+A��RĘ�g����]��r�0v+�5�˳T#�z�W������5�������y8�1?��ZX�#�`���@ ��*i�D[�g��&��n�;_�o|[��@�3�P;Tp�@n�a�ӊa�����6�n��;�1���*~g��M����J��R.;��xrv�V����A���I@n[e�G$S�7!�J�,�E˿I�~{j�ֹ/m��c�78F�xsGj>�Kq-��9���h���l��[��TzN/+=��q8���rz,j b��m� M����&�WBP韺�9[��2)��&g����"(��[��Uq���E���g���DH!Fl��ch�r+\�(?~�`�<�6���؜MS�$a�.�בՄR@�еI� 	A(����t�����G(�V��
����5��I��:�N��<���bϞt���{Ԙ�e�6�Lil�¹�!�ѰrWBj#����
��I��Qjkb��f�&k~�ڍ�E*aL����A��>N�g7��+�4���2�[� ��@àI�j�+N��Ec��jS�yB��e�A5�"�.�*�k
(H��j��їB�;�����m�����Ij��y�Fٯ�Q�t�)��f��{�F�i,T�"z�0�tS�H�	�ȉ�4�'��v5���ި�2��a�������F�e���B�Sϱtr$�f��k����Ӻz�#��h\�1p]s~�6���f��(��U�?sM�����Ν� ��)�3Ћ��c���6��"�������
݅�.��tǧ=�;���+����7
`JkY`t���^�������c�UK�>��uۿ� ស���l�r�X�7���%�J�4p��k>�0�Sp��c��li���Rs�U�)����,$]5�1�0��:�F�W|������H�,��̿>I�9ܤҮ���N
����)�\���ǻ��^꼆&qz�^5ܽ�iem9QZ
�D��a:�~��JY����ʶ�n�ه:90h-Uĝ���*#���Dh�+��U�8&p��:��ώ��P�������I.;�x��4��ׅ��k��yC��J{�T�uF3�Ys4K����2%��I�K��R\m���a�3�'d�V��� �U�b����"I���cXݻ��3Y){�{ށ-��������������xv{/���w5�?.b֠��N����d�����Ǧ籌��'���K!��X�MN(� ��p��JkI��f�����&+��zp	����Qq~o>��ٺA7�ۊu���y>�<-�b��BMĽ���y��D�i����Q���k)��H�%B;EE`앰��V���w����8.�vaݖ?`�IP'�s7�l�cwM[0�W%����ԍ�c^�����Z�r�@Ԝ�ğӵ0���	G��,>�`y��%��xN/�.WK��f6�Jr�4};e&J�D����i���5_��:�Մ>y���P����H�ʴ�Ͳ�t�����z���P"�n4=c�Q�t�}��r�\�XpF�*!Ss~l�����S�m{�x��|­.k��EY�gi�kw�.\��Ln��I����' qE��������r
�1JC^��O�ǫW�%��$1�=�� ȏ�I mj���m�F=]w��_u�p_mDH�.e8.H�A�D����Xx�aF��8�����U��"���)J�&K]�ﰡ���_��Q� �)n���)��X `��(�+�ֹ��<������� xpb,��S�@����$�p	o�o3x��� <+�b�h��P빢�S��d@2�lm3g"ۍ���q�v�� ��� F���CN��C[#�~�1�|��ǅ7�N��� �²�;Ef�$u�M�mE�#8�XG\�M]�)!����ȁ����l�F��ڇ�I^;�}�i71n�p�.����q�J�CQlw�F����L�ě��x���L�%�f@3р�3k
A�E�9)����Vb�^s���n�����/�Krf�m���=���W����u�ʉ�~�{s�1nt�Ʀ�~�D[c��j����ý�Y
���O���i"�@���E2V*�h��i����Q����6ym�;���"���5���"����h�ȳ�a%�H_Wa�v�����IZ����2�Gҕ̉�b�ď*�[�I��%c�5���EA�|���?�}H[���
T��O�����b�L�$NY��	,$�����U~�E��ͷ�h���QOęDܫoۤf4S��T����K�@�B��F�����$.d�W��<�S(���Fqݿ�SI�@�v뙇�
�n�w!�R^<L)�A]P~M/p+��C��^�]<}#�fg7�#ZM��_n�<6�y��NR�3��$7�t��N�/l�z7V+�og�S$�(,n.���$���1��.`~Mn��+�:���n`��/��<7+(��ZB�va1�7��t�[��#�lzG�Чإ����)�ȑ}Ÿ��F0���{�T6��*��T]HP�(�ѫ���g��!.��V���hb���8�0��4�/�{� =�����g�"	l$����Hn�y�~F�e��a��>Q����?&�N&Oq=�膘r`Y{8=�g���Q��D�8�ڻ�q�/q�X9q���֍��M�oQ1(�Ѣ�1�*���l�z�����Ev,~�M1rx�o�������ae��:w�͘��ɰ��5��c�bM]��͝{���[�*��� �X����߿�<a����'@�$K?��b�ͪ$�k�|������B]t�Ѧ��e��5|�<���X��*�������썯Q�S��h%�K�!�T��	e,���u��ܗ���O��>#p�
5I���֐�k�Jr�,;͚���g"��kHK�Qr�������֎Z��K��q垸w�.�� �O��6���n6���[�#5gH�:�<�?�Wx��F�Q�K��tF�mn�(eW�)G��i-���V�8aJ3���ww0e�E�9NLw�Ϥ���w�39�h�܌<w7VEW��h�D��d��Xd'=D��`�+�e�'�� �V>9��Gf�5O0��yq־0�Ʋe1RĆs��"��	��^��I�A"ZJ��E�hN��,;1��q=Hڇu�4R���S�Tac�Ou����$����*3a�֤��}��%r�	F���BU��PW���Ů!��o
�n�fPa[�5 �{,�}�♼ 0�l��`����a�Ak�T���7+C���)CP2��Xw�� �4��#~�F��Ύ��r�Ri5ץ�铠��H��,�d1W����e����O�'����g�k��g��m+f4��ޑ"|�m.�'����s�'Cb��;l�{XO�D�)R��2ِbd��W���j��9� C�B�^8kW�d��:�]	Bg.Z�T�I%&w$�T.����3�e
v>cQ "^Y����,�;�70���A
¡�d�觉�z ������*��Ox��w�Z,�K��3[�&�bJ0�|���N���I�Re�Z��D|��K��=aYu|�^dQAVb&?'�rR��u�KОu*G	���h!%er�K[9_���?㘎>Ԍز���Z1gK����I�N+w��?���k�P��c���|y�Z�#����'o�v=�5.�v��� v[��!@e����:B����Jo��fqI%�&U�� �_��ۿܰ���Y�~�0Xk)�s+����fm��°4
�����6F����!нE՞v&=��̪��P衹8)a>�!��^�'�Q=I������NyG�T
�Э�� �V#�~	wx���A����2��%տ������-̠��= ��0i*UOe����1�;���9��q��яb%M��9��6��\]$�����ZW�������i�<�l���}�Ҋ艦:���ż� ۛ��N�bK�Z���b�x�Qn�a.Х�A�g�R�G!M�I�ӟn��n&~�<���J��X����P<c��I��@_vCSܚ��Hd����\��V�����§���C�(½�������؀{a�EI�1y��g�O�����Gp
���0��bU�/��,V��|7���)2]��]�D���_����:Iv)��jצ�	ś'j�&�ĳ�;AtH�C�Sbw:{܊<]1S_�����ᖖ����,=Ro�z�$�w�RA��'���;n�Xy�Bu�F�8�r�s�����_�7\�SϪS�a��GU���ZZ
�B����~���9�M�B@#����sW?�'�e�ڠY���"1��Z��^��T��~���ęc�]CL��C1Hm�D�	�d���7@<]��)A��֬�lK x/Qj29ݟ���	��'���-��z�:rt]2Kn�</����L
1`��o��|�CG�
;G��[�2q��/LMbL ⧉/��<�MrgJ��yO7�/��5O�U���Q-�Ѩ��T�+p��h񑾰�^�I�ʀ23�p6�I��:@�q��ž����(R����s�����f��L�J:�*f�vX��~�ʄ1�|��]�6"�~o��
�v��lC�;SbRތ&K�oNK;�ZfkFb���#0�_x�b�#1��Req�"f@���r~��{w�O�[Uy��ĺ;��V��ax���d.e�oSˉ������)����oVU�z#��g��H���j��P�XN��wJ]M ��fACņ@�K[�S�0F�-�uX%�OZ\%�wZ얼3M�2:�[�-5���b�3-��j���.L��o�2��}���Gٛ��o%�CE�������z�UC=`��:��I~R?l]����_�{B���]C�3�&i�,&QdhZ�6a��!�`^��=E&9@H�q�jA���ޏP����#����j�o)U����C��9��y�c/#^��/�VI�XԮ2'v�i9?'	�,�����>E�|�Y�I��]�XU�{��l���l�L]�J�jȓ/[ T7��$��+�؟��՟�E;k����8�?�>h_�#:���Y�_�P��O&�^���Ŗ\��SYlͳy�Rh�,#��8k7H~�o�h���eT��m�CV�0F`�̉G��15����$�n�|<��T��[:�q;��n�\0se�=��*���o�<�����R-"�>�T;�@�em&��%`��@G����&��5� YO���-��<��э��gZ\���x����j		�|����ܤ���i���_�RcP�eD �I�#'���-I���܁,�����?`�2����}_9������ ,�(x���nez�`��q�gFq)T��̜=������i�x���5�͚�5�7'>�����z� XX4P�k&x�� r����dF��z���
��j����HT�|^`�3��6ЍF�}Q>c(��.���Y�9.O-Jm�{�B�Ci�-~>���%�� /��O�+���1U,�_��~%�ݞ��&XA��N����5�oy0(�Q�N�T�b�]�I���(������9�$�����(~�\H�聇*��Y>�y�j��SG?�6Dm
��Ȣ#��C�d��`sHi���>dmH�1�i
���[njB�U4�����q�I�F	#1FS���t�]��M�З'���U���Rlζ�q����m6�V�ΚN}p������n��CXz<��~3�����f�9�0%��q�ֹa���������nedҚ�f�_:�ޔHl6�@?��գ3�^DW�V��#�;�L�7��+�}����?�2��3u͒pЬ�u��Drr�sI}�F�d��h8�qh����v�̐AS_��t�7��|����nC���ǳ�A�	 �M6��x�Ǆ$��ԃ����jܟ\xk���I:D�r���n&|n�[���w�uhxep�͞���\���u�t_J� nxD�k�߿ϗ�v��~?s�ֹŕ!&�?���"��,yL��bGЗ�,;��@��`B-m3�[>e�P>{�Lkծ��V��[V��TW�_�D���8.5����d(���3���~� UDz����[�r�e$�=]@�j�,�̘F��Զ�#��@f��aÊ�4�Fm��KM� ������Aa9����r5N2���K'q	Rdͤ���y�.Y\�f]~Uw[�.��}\���O	)0��;�Z>eV�z�#E���4=f���}���q�2���E��tO�����mN����:`ȓ��*o�;�R��3�Pp>�ldg2��S��>�����
ӈ�m���{*к���-g�u�'>Y;O����}`a�u�N�V�J���u<V´���ɪp���\
ǂ�ur�Ԟj/^#�W�M� vb(1����֜�-�À�=Vj���I<}��j]$�(�%���@[xG+����7��eM�D�KD=:��w�"�<^��\\��� �j�|Ը�z�|)ktw��5�%G�~}#2h)�͋���w�F a�?,���F���]����mK���K�Ϸ4$�s�Cݥ�V?�pw�nFq�t�Y�j����� ��o�\@K�g8��$M���d]�@S���{����/�#Z_I߾!�e����%��w���@23��5���(qC֞��|dXP���P��0��fS���JbN��:��&Ly�!?*�5åZ�����7BE}w�P�����7K����=zC���q�[�������Gl>L)���C�!�!8�a��`�f�R��n����2��e�lzVϠ�J���]� ����:@�b��o�K.sg�J�pv¶���g�I��]�+����/��&���?�V��`�����BG�&}��9��@�]cn��"&��- �/��6O��F� �hɠ���s �8p��9�Y_��Y͛H�1��(��:x��`')Fh����&�imh�q���M3���G}�A�]�۲s��?���פ�T�K�J�x�Ud4]�Ԝ��F���@O|���>��n	vm�r�p��6���a"���+~�<�둖(^���FS:U���/^����
��O���1^��j�T23�=d����u}b�qQ��]��m�l Uh�/n�_V"�J\W�Z�Exg;�UdE�[8;�Ib�|� $<�t~RG7�"�� �V�WL��f���,g�WwH���z�z0ӑ���{գQ@������ k��_%���*V
���9�:�� z�iD=B#RE����/���6�ܒ�t��f.;�鲌�?*dT?�#���i��E�[k|��%��RG��2����i��9S	�P�_
��[�A��V�tQ�z��踊������d�U�h����8h�|��x����^D,��Vl����=��L�(e��3WhKQ�;;�c�L��*\�'���Jw�$)��-��_ڷ���w%k�g���ښ	{��|`}���L��-I�}á��9���d������8r�*��Җ�ݐ��)���DA�
�	O�#'��I&�s�ޝ��c���p7�1�o�$�/ė�E�����ZC�m5v�yW�Ev��/�0��>�E��ٛ���Ԯ��Ր�h̭�4�|bT��I�P��Ė\�t�;|F�x��8�Ԙ��Z��^��vR�����>��K��&�֓��]a�vجo��F���F[f5��C�~�{��"�n�� �uA�����ն��`���`�ה��r���͞Z-D^�IJ�?��H����ݺlŵ[�X����yO�*z/��kԙ����o��[��tI�dṉ�?�y��ґ��\e��
.�g�/k����*`Z.PF �§_���0gI�U����l� ���J��EU!d�+C�}�� 
4(W�~���~۶ ����RH6Εm�����
M��[�[d?ȁA�yT�\R¨�+]'#��h �2���-�aΞС���Cǹr��b#�R��xd�����������ÀD�v�J�1�U��X��N
�2�۫�4熐����X�[	��?�q=���lXP'��d���>_Gȍ��/��w��0�DShbb?����>�5��v���V@�g�W�5v�l��%��rn��-�dϗ D�`L3��waF��!�oS�����Ӱ'!M��&�a=�$����#P("p�&����Y ���6�mt{9(܈3a��(Ae�뉼#^�b㟤����h�� �mdrόH��LJ��F�њ;��5�<��?������ի�������1`}F�X&{��aB�8�`	^��_�j��]�����ɸ��?����\'P� ��b��H�E�bu���&�d�؟��E�Ϲ�������FVn^�c�5T��3px!*��
VT�S��mќ���7�m�8�JTm�ܾ������2��r,�-�ZcB�BB�:�S����V�?�&eVR [�R������=�2��L@������Ovo9�Kz������~�Ns�������#��c��sŹ�ߪ�4�(g᮰YL��K3gC������SD��E;�6����G�!��:!��Bn�o�R�,�1�Uo�{�$�8He��dsN��؜�,ǢUy���z�t�����o�],��VOF>1��%��H�������ۚ��_�y�<�{�\IQ���)KE�-��;(n̗F��"b�-#��N
�󉍸�%rWlp�l?0{���L��6�o�M[Y� &y����	�  �+Z}�����<��jH������j]RG��=_�����V\�wsr������!"j8*{@&~Hf���v6�Egt.��r]�<l�};�CP��M��i�K��t�u���ND�@��5�r�~�N�z�aZ(�)Rz��(B�m�^'S4@G�^�0,{Uo���K�y��ҵ�a��I�d�+�vb�
���o
2±�O��L�v�Q���O�Y-�:�no��s���n�|�r�p�RV��2���Hu��&���TΞ���,��D��d���d�f��t�,[w�'&��;L�.�{��1�Ф4��'aJM���|�G��!j��͊lƬ�aΕ�c��I��`c.�1���)����ն��uC���b�Cq�� �!�]��F�jr����1:	���& �JMFu@*����m���Ǉ����= 1��� ��ʓ�M)/$1�Eg��J�BC���k��Ix�����3ȇSX|.@~{�)Gh�U�s��l�(��|�kֺ��D�^���`�����#�O�"qV-aN�ne<�7�p�a�)Ҕ�",φ@t��9���Ýs���Y1��H�>�H	@�#{n���C�>~V��$��d����ٌe��Yn4e�����a�q�Z��@��{|�o�"�Ӏ0gƝ�.��a�5ɛnGz���bQ���õsF�UG���Eκ�++�X�����Wm�7�U�&R�r,Y���|��i���9j\��L���(4���?�ģ2$�":�fD9V/�z���U�O�+��W����Xфʰ�0��#[�;s3���ɗ +J�]\��m]���A\��q'� /�U�Z � Z��r<�6rI�gY��j����
�Ə��4�E�[�WCs3�y��nB��8��yZG���+�/�W�ҦE{��Z<C��7�ƐF������'���p�1��`b.΍ˋ4��]��֟��W  �a]�ˤjD`ڮ��k����\h��|���D�!���p,(��S$dܜn$���ф֣'��~��2g�(��ը��9��-*�I'�'��1�7ę��y��{�I`i(v?����4j��Aڭ��Q!�R�n2��=#������Jf+�������8@���q\��^��Ơ����
J�lq:��EX(G�C[���I����ɋ�,|1�"�uXv����fj��9�b-Q�!�#CB"�)�4U���%���f{�����:"d������n��UN�ݪ�6vI��XC����VP�2 #AH�9�DK�f���'>��7}ע�S8=z\BI�0"�oșm�P�;�So�A�ߤ�}�oz@��8& �Nz��5�:t��,��a�N<��ߢ,v�kϘ��]o(�;.���s���B���@~8��$����3R�.��"�q����S��;Br@�w��J��8vY~2|����A[ /�q�p�;~Z���X�&~:��ۏ�<}1����Z��P��,¸��~�(M���XnY��Ea�et9�ƃv�"�Qh���Z��^�~*(+䵸#�-�޺��t����-%�V|fLg���vF ����
�G�vK@����4�.�DbV����ׂ�� ��Y	ω^�Z�?[K�BsQk 2 ��Ѧc�+}Y/Z�I�8��,�Ѐ4��q|�!	^�q����2���c���i(����Cf7�B�ͭ�F����m>��=��9���ߧy��1< �KE�h��VP�p[JFm�ش>nL�)0�p�E3{C���Mu4{9�ʃ�p�
A�hO���e+&7.{��#e֜�嵣��4�1�J��a���[Z"����������"`��Ɗ����7\�E9�1����|D��,�WM	Q�� �b�菦|���F�N������Q��5k388����̚_�!_r�Oad��ï���Q��k����[Ȟvҿv��
7���A]����4#l��#��-&��@|�ƥ&�TϸE�1zz_���vr��~5�p���g�����ҹxѻr�ֵ!4���ʫx���>���}�����S�OwE!k.G�^J�
.r$pH#N>���!I���ѧs��K�2a���k�Sͫp�`UPas{n���o�u:M�����-HD&� :¡��j+������˿:)�v>nZ�
�Ed����".{�^g�aT��%⩔e{�����F?�15��'c7qJ+���?�ױ���e}Q%s]�����
O՚�v� *��
Q�v!D�$��i4`�����r�ǡ�8�>�	F'�|����j������]|n	ˁ�׵��z�#݌�g�)C�>c|����L�]�l�Z�����o��"H�z*/E��#�B�˗I���UE�Z��Ի�^�C.0�@'��aβ�����|0�q���4�D��f`�.��M���n�LG��M�kHy&x���0�h�(�����U�~#2�����h�!1"���(E��]=����_}��M�(�pG�vg���56�̱����,��I�z宆��`��=X��l���'�AO?��j�p��	e�{koI��!�>7�Πy��~&i��6(У���$.偼���տn����)QS���3l]C�1���뽀Y�=Ԓ���54���S)�q�[Jp�2��[��\n���z���;�m�o0��_� cT
�{��2-um7��}��{�ɐ��Y����U:N�|�!���@�����c�A�|�S����bg�h�D������xlLo0�`/��V�^v��֘Ĥn��١���C��6�e31�+b$e(�Rr5�:MY�d�!X����$Tl�bX&*�KY]�L��	3�)	Q�ߒќD� �7�=�^�
�VR=�B\�h0ç��K�<��Ҫ���h�IYT*��`�М�����9H��1CX��3��GH�\c1�O��I@��qk�����xF7����Y�����}:{:�L,�=��
7q�C�!�c̻rS�:�L�$+B��w4�t�|&RyOy��P,�S��k�����V�C'�?ܯ3��8��x�IP�dP���z�D����/�F�f�"����-q�/��_���0���4�B��a~@�<\�[��B�����e{g���6�7I��_uU��/��p��*�������}� D����Y����$;#�d�z��Hx�*o�}����1�o-�y��`jձiH���]��]�J',�h��!
��jz[ �����2�ތѪ�%���b6,}�٢_B�y's�M�9FZ��։ޝI���8J^��Τ��!�gص6ˮ�J�aӘ�h)P���N�˽�?v��hy�^(��x�}b����
yt�2��]Ŝ뺽�� ��i�*d�5�+�� LQ�ʌ~������2�K��=.1�o�1Ow	:�~�64�C,<���H/��buY���h�}|
]g^������9�g`��p��b��r�ǰ@!�������bM|�u~,��=w��mVC�i]u���P��? o���s��+�*��v� y�.}ƀĸ7�8��i&���(�qR�Э_4�?EU^��z���;�7�}�pa��Z���b6��V�w|�Q���q{��+���1%��
��0MW���M��1�$����MZ��a�k���o���m��^N�M��:{s�պ�"W��Ӫ��V8Dv8ip:�U_Z{)7M�]�J�z����g0��)��2&[���"���P��=I���-�]	!�i_6�8�=z����5d�Z�x+�7������3����!��st���'�7џȗ�*ʘJ q)O��)�Y�w�a��Ǆ��FE�V��q�{@X2���Z���N���Dֽa{kR�K*D�L���s}i���7c.�g@��P�Ԉ�gԐ���Ӽ�`\qn�0nO���0K�R��6I��|���E�h��b�{�U�Y�������G��I��"V&~̄ic�ʘJM���#�Ӣ$r�������6o8�+��&��D2^ط�ټ��Lқ,�z��;G��g�뾗��;lȈ��E�Hf���G���w����v(d�{��G_[���j�9�ёm��x�<ҴL7Z��9W��:��x��ߴ��AD�+�@x�Մo�Y	����r#�ƧY�d塒��\�b`��e�}��*��,�,}\��$��I.f}�7蒐C�� `ı3�ɭ���m����U.n��=��t� �������w&�����0NPp˩���$�Q�8��+������bSiV��*/�
|��W,X����MR�Wg!ɺ�YA�p��m>j�`�V-'@= 3h���)�M���
o;o��]M�����������1���y��BU��r
��+�*�KN �z����e�g=�Z�Q��ʧ���B,��D�x�-��l�LQU�fb �&oˉ^;9�~�Ŗ_�	���]'��д�ߊԪ����YPgj~�$D���, ]h&3W1��ptS8ig���y66U�u�ČGή�G)�^�Y���E�]R��fN.';�8�?)G��V���-_n#N���'C Q�o�h�c�t"��?���pGI,���a
3Qc�G:�sH���GT��=���&�����ʩ�"����10�f�\9;Y\"9�r�p/+��XC�̻K����m�J'"��߳G�m4�7��0/�[��7^��4���U�X����'�1\A�IG�^�L�k��C��]_;���\t�!��\ZU�(|U8��_m� ��%�b�	��;K1��g W+L��z 
�:�~��<0�M��nvee�&N%�r�4��"����-.*���A,�}0y*tF�ްg���]����8�5� ͱ�=�%/��fs��P�u�%�A������.����a��α��"u47he�%U0���P��,��u �/��#��t���گ�G��^��Y�y'�&����#E�q��ۇ���f���f�e �o�}��H�U�B�S���'"frM/ ���Bǚ5��6'�%Xy+�sUm���='�p���(�7��Z|^ߦ�i6 ��=�
�B]W�O�s =.^p�&�0w~hv�S4|ɞ���f�(�ǀ��p�O5@TxT�	kU/&X�kx��5ٽx�<�^!�_�{����IŽ����5i���h޹+KfD��a���0�+/"�nÆê��+M�C!sS�� �Z�&̔#=�zv��P�^ji5�A+X!�yc����`�D�ʋv�z�y������ 6-	!i�x~@w��]��ps`9}X��P�dpk��P�!��#y+��[���]��g��_�ό�b��c2��K��\IT��kR	�P7!قל"
߷�]���W�U3s�P�kE�,����/Ժ�_�</s���@�m��)�W��ZZ��F"[U�%M�H��NңOP�*Q�K޵k�]t���\Ե3�!���z�=��M&���(��C��)z�K'UC���4��$�7���櫲���>�OMғyP6��s!��(��w���ER��K 5�D��ap���l�o��tM������J�+�Xq�/��ߤ�Ic�鑎�"��kі*�s��%Oς.>&U)˃q��y͈�`I�A�`P�^���Z����!�����l2�~K]�/���-on@``���2�@��"����$��T(tb�Fc}Q�i����h��M$��w�z,u^��(47�Md��-�2,]�����K!��1�˪=J� �V�k����jڙ����ꄁzl�A?m��e�t�Rww�fs�zj�zi�l�WQ����R�l�T^��P���-�6>��� �l�#��Ba�~R7���U��u�O7���F�v{���31��F5��,t�6�`ԟ��4!�t*{�d��^��޻�A O,�����=U5�ŚX�6�@Ť����g����Mp�������*"�uH��f�F5Н
O��7�/��INz��A��8��̉��ۅ�k5A/�"��M�s_�Z�v�cN.��<K�����[��HV{L��Y�q�F� ̐�:~O��Q�@�V;�Z�C�y&��Y�4\�3�myezD��1�._c~sϫ��:��M�e��	u�{�AS������{�!��^9����3�Щ	���EX0����'S6ys�����-!���jo���5�ɟ짱oY�R7w�<�Ya'rC���&�Y�f���	:�����	����{L`��&_�ө����%9Y�v��~�����`���(Vδ���	m�����~��Yg4�W���B	�@m��gHm��i�0�s�ǹ(�����G-�2�ў)�K]�����W/t
1$��c$����PЎCbv킷���f+,��Wi8sl~ت$ٽ�[ou/���fg��`9�
��ff�s!��YB�ǯ�w��͓_�H��]<P����oz�l���1qZ�]�;�X��DV <�zs��0@]�F酜[١�=���l���z�Z|C��y�km�~�����3�Yn�4x��6?�:2�9�z�
��Hė�ߠ�A�,��jY�Y����N�����?y���d,����⒦)�%څZdމ�����v���/Nݷ4?�^5��J 6�Oc�L��Gf��R�p�Oue��$t?��=���_�	m���>Ĭrv����R�3�B�SLL�0�3�w%_�� 3�b�Mj�bY�d]-��a����}���c����͚���NK;���P8@�a��*��&?c҈F\�!�с�gL�%6l����q��NÒ��w��40b�A<	�	e������V댡�� �<��	�Ek�^MR����$ue��0�b��П�Ǿ*����=3�,�Ye�Ԧ���3���Ϣ��ZxO�8+8L�5�_�
�3�%��=��x�#���8���=��<D���@KK�ȍʃ��?�H�;��,q�O%�ȥ$K�L�_�7�=+�h?�S/e��q���q?l�ţl�/�ʻc��y����
j���}�Q�h��"ཟ��e�?zD���=�u�Z���U]V��7!MDqLj�処�LǲR� �hz<+�G��&����(���S�QL��ի�ʇ�����(��h�'V�P]�-i:eG��*i|��]Oф�W(nc>�©]�hvx�����PZ_1A([h�w�N=��H��/\bU�}�D�ƒq��{�QU�o�ɔ�6ZS끖F<d����6�	�i^�[�?�ϰ�@�;���&{��>#"��4�N{%��J��b���v��Rl��#�����
�[�S*�^���١rs�Y6f����١�k��*�� k� �̳���O���o�i`��ν�-�]����*��A��������yp��?x��5��R���(og�Ӎ�8yd�B�7����y1͎?��f:4����Q�[ƫ�"�,{K�Iy�VsC@��є��{��2�f��>Ln���> ��ZpN��F������*��nP$��p�H8�!��T�B�V�$r�H�6�
�j��?^�%���կ��M�0�v\Nv�?5���EUMl`?t�~0����xC�Ӫn,H���ZM%�����k�5%�ۊh����9��:3a�)9�����j��VZk�=f�k| @@ذmð�������9�n���Hc(���4�v�(���#M�4[vKZ�~��NE(�z�D���T�^���^��so��[��;���"�|�Qj~-8ZW%��N���XX|^����`W�w�4\�x�mԺ�I[Us� ���{H�	c��q��?R`�wՙ��A
�m���V��y�&���?��	�ƃ|-Φ0>W�2 vC�uD�����E�_�k݋�ɿ
c�J�����<��L%�Y��e�ӛ_��a�->.�tP� ?�����q�Tʷ,�F$q��9��u
Z�x�;�̞�A8�LxF{19zIN/*�pD*�^L2��mzH3>��mL�����u���Ǫl"��V�9�+L⶗jA������5\�p��4F��c{��F�P�\C�C�M957�4A�����J�y�'LLQ��|z���a<o�	�CLO�s����p����k�3�C��Gg���s�.�姵��ax�G*�|?մ�NHڿ�c	��F�P��d�J�MF$�]o�YO��oj�"�6����ҾTU��	9���;�>���FӢE8��/9mT8���9�u?^�+�~�aG�",�Exބ�l
S�h%����8�	U�%FR0�@D�gb�O\d������`a��}�.��\�ؖ�*�9��q���Λ\����p�;�V�%*�m�Ph�nS�"��)�k_����#���5�vn�gC8![OÀ*�܄!D��WN�][�~��>�X�e��"�������q�:��ɼ9��m�R:�K��T&�F�f�:$�>2[땫�O#���N�S[�+��)��%Qh6"_y&B����!��a��0�.�c
�(�5���'���U`W�,��w�8�����.*l�v9/"nx8�5�Z� ��x�����U�a�@��;u�e�-����}�>"�P[���3�Vl�G�w�u���%�ɪ7��K�/�aX���Q��=(Г�?��m��f$M���(�6�� �
��}���:��::��儈�auB��ZS	��b��K))@	嬳��{�ϯV�.�h]SQ:zo�_��{��V?��x��êw��(��%(n�Kh��k1��u ]���G��)����e�vH��b����U�A�Hg���#�+�<b��(�ݜ��7�S"bXIm5�B{�ǑA��Fu=�QI���SO_�ڏ2	��������u���9�v��u����$3�{�A�	�o�-��	�'�����U�3N�J���~ P�$��'�J�H���;Ge��o,���&_*� ���ض�,�<�[��]�mF�wM�ߪ�U�}9M��f���U��A/z�)3��J?�y�P[��]'��>#��Vw�+��\({�pU]��Io��y� Hn('<��$*,w� �E	�md)b�^���S*���h�M���n�2��h��Xd�/-���cK���0�I�
�6}z<b���˴n��:�a�����=�O)ZC�x��@w�̆#6V�E%2U ��Da}�L��&�<�<TT)��j�x�%e+Be!檐b%l|���3�	��82��痲����kq|5�����4{�u<����v3��W�N3ksӒ��g)�����W�k~�����S�e��KO��rT��0�����!����wBɊBXV�����P"���-�x�Iiٱ"C&"My�	 �f�mK�g��EL����R ���+�F[[VC�5��ܳ�f��Mr�A�KJ$?�DU�n�v!}!?9�*�#��/���M����@� ������P��rSFX�7iCe-"R�9�ཟ�r������w�d���k��Z��D f�!�J�h�� �U���A.�,R%d��ޡ�<��O�b]��|�VVf� kg�ֺ�m��txۛM(���k"UPx����6�F(�M;P��w�q�R��X���i��I�4�?

��d������=��1�pIUX��� ��
gu�J�!���m�r�F�^X3�!.�����j':.[`_3m�����obs����6�����S�����d�0�<H\�������^[G�/���<9f7��Ƈ�6�h��y����E��a_g�yb�T��%�G	)=)=6�����F�B-"�4sA>��QAL��:���$lrP�{�2�3A�ҟ��S��M^^�������H�= ��센&�U����l�w�d��"�����\t�-i����&D�ʔ��,3z�L0����I��s8P�ՐW�X"��uz���Y���S��ڑ��v�[�d(J+7Ԅ%K�@08�¼h'An�8X]M7Y�$����;D{����ٽ�ZC�}�(k�����
��Ox�)S��P&�1^�������KS�ӳ���$0���oF��}l2oi���N�W��d^bPd+A,�z��xv�YJ6aҫ��ߢS������Q}�oěA��)���ɽ#�Ȍ	����x��h�(q�Ez���TR��e䗼��t�H� E��D���F��W���<���ŧ��E;K�(Z �T����X�����d�o� n�{���,��@�ɝߞi ]�='b���Ōk�n��.xL_}��M�o�#�_���W��,�+>���!/��Rv�����	O�ԝ֧��g�\5���#)�rK^n
<�9�1���Vv#'zT)U/Y� OfT�C��A�RUs��<r��ګ,E�9Z�&O�2��u���^��Y�Y�mc���@g��2�X%��n���X]ط�"��,lC�r�:��}Sx� ����Q��X*�We�d�o~�Ln�8NKL� f,$n�g\s�g�����G��h�������R�[0Xj_��rk��ct�R5b�!Ss���K&���XF/�����mW�֋ߓ{�[�?UOIx�[\,��fqo�_��'<~^��qӳY�L{=)�la�9#�@2��E��3[����y��D��v�aW��Č�/����:�$`0����#����P�83�>#��~�p�s��%r�Uq5�V)���[B^��Mbc��O�}M���� ��l��� �����4��f'#v8q�u�ͦҟ�l�<����R#ӯ�S������,ّE��X������{��ajD�]f��V̢����
l�K�M���,����]��~4v�N
|@SV������s��+E����eM/ЋNU��3��u��MIC��CQ:�6w��0H-� � M�i��%��DEG͗�<������ht�>�0J�sO��	��f��X�Ss�X��c�>YF�gN1��_ę��Ff��r�M���q1]��c%#��E"��/�{�T�a�8���y�b���mv�D���D�v�����cqf��T�����e��MBٶ�5W��A�w�)��U{
��q-�=�hZ��&��>i3'aG�nY8�L���:լe}��0�=Kն5]��q�a�o��_���g4x��n��}α}�=���[���!�)Z}K�J�}����BL�`��x��K �e겠U�i?�ۥ��41��0���:s��xC�	ƚ�>q��'*��s���/�
=��S4e��c�������G�ƚ�il8�l���It�K�I�����@��μ�(�g#���4��6�ꍁT��G��z5ϳ�*fcUnTo�a{��)XU�y�hڜ&Z�����uc��F��h�P�*���b�EO�^s�Vπԗ?��`dk�C��w�f�Û�E�1�#g�n��f��G��1�W���<͙=_Η�Q�>��/��v=� �l��\�8�����f�����Nrj����3�<�;�g�2Q�a5�%|]v�����-�)��t�^�P��ݨ��s���{Jj8i�����c�2�"�5��(_��&� �-��� ��4��f$�xu���bx���8��,:R�Z&�G��:7]t������;92�z�8�Un融�+���d[yq�*��\�~�ޑ�&�(��Z���shL�G���x�;� ��_��{z�/Xm�>
K���t�20.��jW�^�r���mPYr"jF�=�h�`�l��a:]mt��p������K�)/�����_,?�W�0�t<��B����������[r�56�^?��'*p�O��J�>9��t(ceڹ��H�}��zd�)3T#�jwd��H����!�:����Ŕ�p�o���4G�aÜo/rH�I���a��tc&8�o�l3mV�O��g��w�DNi'!�1���5�,E�ϝ��'��+q�\�WJga`��ݹ)7Y��~2�9C���ֆ�o�R���xwm�]=q�s�5�����G�sC
�V��E_o
�����{@�j�勜?�����  �ٽ��t��m�
��_���\�J�O���bv��>?�g�l�����"z{�����?	9(�I�m"д�	��
[�pT�u�s��c6Ь�21Ǚ�ӏ�Vr�
���;�7����3���6��C����P���U+��0�5�C�/R[�ô������Ƴc/!Ɩ��]����������(���vdQ�Q��G��n�gŸYb��_���
X:ܑ�1#��)E��t��(��Fe�P�T^ܡ1����ӌq0��jȵ��[�~�d�'7[��&f�Q��A�pŒ���>8	X� �.��F�2�ITf^��%��ږI;k��?�<5���hJ��a~�TJ�5��g��3���P����T$����c�g�TڹW�0R�%�T{Wʦ��j3B���mF�^�<�����k�j�}���q,��q^��K���L��#��ݠI4ii��M*0ʔ5^I=�ʔ�il��y�rV�/ܤ+=��c�F�v��m;�I�E����:�����)��!%����k�%5�"�D��kL��~���6�M�:��T�p4���;l��a@uV�� 
�H/s�r�K��G�,k{���u�(�d[m.�(�d)�i��y����D\
W��A-��9��_?SM���*�)U�)y\�ݩ}Mo�p�R�X�Ѧ�~��D?ҵ�̣����O�J�p�0R�M�v'M,�pv]��^�����v��;����0��aj}�G>ޑN�]x�*H+*�.��w��oc"�K��<�5ލ��p�tW�vB{pf�0
V^��tC��<,������ȄU�(�]1M85��-�8�A��U�E���n� 5m짐!T4N����JG����O�]5nJ�a%*��B�(���c$����{Ѭ����N�� ꮵX��P�O�lQS/�Ys£Z*gTǋ��t-э�
������-�.�N	ʾ�Dl�l�k�u2t�`�&@p��bMq�A���[��8<��=E�-h��=�}Ñ�Y7�CE@�g��I��ԨN�_.z�� ���5l+[!?�bQa��߷�F.��e&��&�y�g6�@�v��F~dx课��o4��oՀF�v����;���W�X�\ⶹ��P �z̮���C��v\�*y�/5s���
���n��	'[\�x�3�?X#���~��2��PD��96I=*Q7�I����ioK�(�.Y�ִ~�j��Gb󆙦K������#����v�"uF���|ԏ�d��4���$��A=�.HB�A,�ߧP�(��!��e��EH������zD�C5S5P�y��4碒w|pF��
P���Okg|���${�܂!� _�	���F�4������|΀#��B�`L<����u�ʥ�ZU�W@���1Ih\3��uީ7�y�tl�����O�r6;" bc�F���0N����g�Pv���?e1�6���J� �F�"'I/A�J�����g6Q#�
K�2]�����T��'f�ߎv, �����!l@,�G#3X�)=Jw�U��l�tݖ+�N�Nt�n�i�tਉ�S�1�h��	�S�+���	� '�i�.6&:��#oc�VLV��g��Z�j��T2+ŶXAV�W�D��p�~��ρ&��Z|Ҏ������_�:E����l�(��J��D !��<H/	$u� ��&��X<��Pq�5�j�B/!s�p�xm��o�^k�Z�%�d�0�Q���J�@`���� � 77l�z�7A��r-��1�{�+�0������B��*�����k^2T�qo��P�7U��`ӷZ��=M��S��ޟ�����A���E���rU��SX�����n�u���d ���)m<�Zf���d�[`�Tv�V���:Ôo�$�F�Wh���bv�Ky��Q۩�j���oc�h��?f��e��S)K����������#�:�f��JzW�	��aj���J+�@����MI��sUB\>Wng6?��}N����C�n�$��*���PX����ꀝK���9?�E�[�3�%�sͧ�a͏X�ζ���s�x�e�,�8Ca~�px��� _��u�W�H�X�G�S�?2�(���E O�pĽ��p��#�Th�F������O��׮D�`�t��lI���sxK�*�L�t1��p�>
ɴ�j���wBPЄ.N�0~5�ȸs��"�|q7��z��ڻɓ�܋�O�����J:�^����P�xiYq_�'�(�j끗�Y&? e5�x!����"��h͠��JB>t���J)�m	f����0�����I�m��H��g
1�M{���� $��tp��^i�w�X����P�|e.2�������<~bhcFӔ�F�g{�?R��v7��J-o?mj��;�/Hd�A+�@ݍ�N���|��b4�S�E���1۵w��>�?��f$D>or�44�$R"1B�fe[9�'�3����)� ;�]ʡ�� �B�
d����޿En_���b�I�<S>��u��me��n������u�/����4�F����!$�6�g��vh�;C�}z�A,�]��9���� ���H��� ���@+?e�H�qc{��1�%��!�E�daVL�jJ�:B�qu��
25��,�<��H���_����������Ge�q�KO�jy  S�U�!Y2�E�wz|�����_JeA��Hq��ʨA��,�Sa~ڣ4�*Uʬll���w�r���R&�ft�4'~r��﫭3��N��/���B3'?	��H�X��_���4{���՗ز��D9Mg<�jNF2�考(�Y���p��7�"� �8A���~+��&�R��7���Z�!��;�Q�P��x_�4��Uc�4[H�a̵e�e��N�\�6�����J%�S��.�[Ǣz�_NP�o �K��e�q�0���7����wgE�%P�, �z�a�֬Н��[<@��r�4�VSd��ڧ8G�. �a|�?M~�� �9�~�
p�+u�3���Ƣp��`
M��$=���~��p�ǅ*�>����Z���xrs9��c���G��U��� ��桝E��SW�hΓ�3e��cAi*^\�β��^�0�I �Y$G�ܻ���+{bzJ&.۰FB0%مr���+.q �ҋG��w%���N}^$7� �a)7i�w�zB$�'� P��88r���a��8�9�'���� ?A��u�m\S�{�{w�L"�O�HoD [�
{��D��7<HS�?��B,|hHg���Ex%hAܤ��(�RC2#��[��G�7������~�Y	"����^�o]�af_k���̇c�q9�/��#\ϫ��C����.�}7
Xr�����h�Q� ���Ԩ�)����<��3k�5��[2l�ʛ�Ҭ����%;"�\�y��K�_�J�uMkB��j���d��PPd�Qݑν�ŉ���Z��\E}��)B���E�=f��*����:��n�
��o��'�������4�x{�:B�fH���#��uߏ��L�8��2]�g#��P%����~sw�SC�9=m�E�]F��������7���&�<n��eћU>��N%�����bz�fCg��$}P֩I 6�tP9��p�������Ե��� �z�O��/.{Bj���N��b4��N�;'�&��m
U�c`g
2�48m�e�x �펥"�N���z:	 ���=�TMy�h+��7�5`��֡�'�Q���;qk�h��,���鼹�5�[�/��d!ڧ̽�5�e���-'=��7�]6t:얠r�0�%T%�=�uoPf^j�dvY���Y���FRg�|b�j(0�������02���g5�������c����/�zO >?�ŗ��<���W���91޶����vR�m�՛t�<����\UP�
,�M9���ix�`A?*��y�F���s��"��et���w�$lLߵ�jX�$Wגl}+�Ҡc���k�����8IQ����+�, ��O��}����cɍ�PQ�g�C"�7��QY�8��&����n�2�?�C�$��� �c3���ɔߊ�0��c �Ҍ�R�O0 C;�1�꬏P��Hew�K���3[(�nP�4W���e4�@tʯ-���N�?x?I�9I;�N��vXZpت�w�3@Vb� �@�\��c.W/i��]�ڰ�0��62�d����y^�pgX�U��bq��Լ���Fe��R lBY)�Z�ޢI�!�yE��F��4ɱ�͘����SV�:&��C�[[�YG��P��%-���<�U�/�,1ʂ�Q�����Xz'A4����
���|����}Q�?�*�����c�� sz$�<�{�<����«��?v~F��<*�e��hH �݄an��m��L�%i߯r{(g@.5�ٞR])�����cN����JC�t��VL"�SǕ^Q%���4 :��4�(�^&���w�ӝ��u:��r)��t��pчċ�X�3Χ?��m"�<'M���Y�/Z#zz���.��'��ɥ���^�=̏������-���͓D�S��s�\��$ʎk�����Uj�k�k��ٿП�k����T��pNY��z�^��6��ͫK�&��8��Y�����'9唅�����hzTBI�0�v/vA�'�'*�n$��um��p0Y�m�?�:{b:�%�
���j�%ǧq*e�ݘ���XjN���}�6e�8����mv�x�U��_�E��I�&G1G ��8�%�ʯ&xO�3����.@d �n)�?;����>��r��e���ӏ*?/����"��<9�ܬ��d�L���������-��Kh�EJ�N�`�z,t1�X`jߪ{��oZ���  ^9��t�Ζ�e�Mq_Tsx���Jx�ظ`�s�Ϩ�YhLX�EI��k�.T̀~0��r(5�9GD��h������銣�bd�&ks�S>��<���4�2}YA�������(>����o��k�޹�� C�����ɏu�f�ZN�؀�� �'a�����sPGi{�	#��<hf�.mKe$oۦ���1ݖ��\�)X��4�Q�A��&��s�t11}� yb��e~D��h������##@�g���=�<��{�@��ȆFD]��Eyz�b->�WD����gK"�+�@�$�(f�v�(��{G���K�C�> �2�>��2�U
��2�䕃7c"Y�f�� � <����^��f�M�W�<Xn���ȯ��bn��\����\��&���7_=��4q;W\3>�[w�gh
L��5�px7�a����:"�9������=V�f�],��v�}י�d�FE-�T�oȇ���7]\���[�r.J�y~UV1<ض�?���A�wv>g��R�˪%��mJ�T�K\�P۷og�X�����hI�4>,5�zt�R���;�����2��&�(�a��q<m␿?BB]۹\��L�>�<�,�P���r�颿{ܹ�#��k]��is�k�� �j8,T]����i��k7��4���[�AP���7�h�.�<�jќ�X},=��x�ྷt�e �¹�(��[��0*�7m���9xH�}y���/�.e7�@@r��_��l~fĂ=Y�~��AL��fyX	3�MlA{�
Dz �A�e$:��c�B�i�)�^YH�`��i[C�]?���	T;M���2�^� �g,-���/^�*��t�./I��Ư��,P1˱yvvw"�)4�*G��BKEq��qjZw�'��n`s����3b���rc��\F�Q��������b2b#v�Q\����ׄ�0�Œ7�1�y��/fҽ2Po@+�H�mLt���9�H�.�H�C�1f�c�����,U���[I����A?��G��� �RaSά�B��LF���ٓ,(t刧'�hG=RF��j�7)XJz4 ?�\���6A��UV��:X%�K�ԥ�L�o�V�L�I7�Ɋ���&_�u�B����3aY+���ty���0|�^c:�K:X��*��=X*�3��U~�6�X�=�����)>�Y5e�h��5��[���ȵ�Ԝ`.���B�܁�Q\_����7&eN��?�ꠂ�ּ����lHD�O�w�Lti�)�q�z;#�1�� ���e�փ$�O��P'%�<�ѱ����Q`tu
a�La��2�N�7뜙W&�ZW���z8��d��E��!a����B��KU<��Y�(��d������jK��KK�w���U
$z+Uc0.�UHӋ<t>9���w���ť�q�{�����c���������s�F�ڪ��v��x�l!��1�c��|�Oe�I��=���d{�K�EV��}��������f�Z�ȣ�昵X�@2[�ZkN���nPn��D������������хJ`Τ�p�r�m��Cy�Tc�#1nS^�q����CL�4e�P�����o���YC��諩���� ���
���<~���Y�l�EG�Jۙ>��j���V��b
6��b_Ě�#��q���ͩ���y��m���w�?}��,z�2���j�P��+a'&*NB`e٭��"B���w, �O�`����:fVe��B`��C���?yX��?y��
�K�����Ԙ찾�)N�0)G�Q7:1��� �5p�B���ע�[#��sS�	6E�>1��1��p��7����|c���QLS$l�k~P�.�b����C�Ɲ�[)���0؍��N7YU/R�~l��	ɒ��t���
9�YߜF�U����|�H�B��Q7�GQ��a�>1L�[�Cܷjާ_9'J������߼���%���4Ȏ�Oyڝ�Щ�PcG-}CǄ0.*�g%w��LgI�1�~�%=���L��F�n T��{@����s���8����������h�> ���K^�G�'��gh��ପ��3;l�JH7��B�7Un?Z�ʬN���82����k;+�����N��jK$3�(H���x��p������;��*#�<c1���~��wU�"�W/2����g��w|�IC�� ��e�c0�,����ե��<Wi�C�����=��|`4��G�w���,�t{�
�� r�����R�yХ��$�M���lM�Kb��pN����8��g��K"X���Yq+h!�*o	Zs\�V:"?�`����1��|L�Ȕ�p~7-C��y�0&:ݔr�j�Y-�)�h�C�Nu�ƙ�F���{j�I��w&��-�	>�@��f��_�^{�����k�En�1��m����/�)�LR�Stә.ZVi���˟��^�m⼑����d�QF��(�#y�1R�+F���h=�;�L>&�"������!����m��T�©	�7�o���L;�d_GM�B}��<�8&�?�C���?�.�����&�M��OS�%n]&�C��d��DI�{�E��l�
9f�a-A-���0���0YE���|;��ҋ��������cBA���s@�~��L]�j��k~�r�r��V���C�<:Ur�<x֝�B�8b��|��k9)���Z̉*�����5~��=oi@��p>�m���S�A�<(�zC��`�W�5����[͎�t.b�fS��'��,���%�l�Ժ��o��׺6��|l�︔�4�=:-��ځi��]�����}\�Ce���z����b� ��Z�3��� ]�������L���sH�
Ԙ$�ʰ�N�D��� y�a���Hd���E~�JT�,�t	�h��V��b�a�I�bRG��L����1lp�0|`�0�&@�����Yb��j1��?�Up���lbc8n!2��]�^�C#�˔�;�C�%�Ε���E%v.�˴��#n²��=kUZq+�S�$���q�V*�X��Q
3y�>m��A�_"8;��KT�Q��$֬l�c�Tս:h����e8Fbԉ,$Ǳ9�y�Ŏ.}�<�*(D ����m1&��7}�.�{�:��('�%�T�v2���?��\-Z�ę�q���k��QpԮK��AXFy��ڈ�d�a9���n�;��,�U�a8�L�גtO���r`�NX����h�ߠ���̘OJ�s?W����-����Sي��`
��Ơ����[x3r!��n��ީ�⃺�bҡ7b�v9�\�(������d�M�t�+$�׹1a��gcD3S�h��R��gI�aK�d/N����o��4��-��C���ٜ-P��E�B��1���:��
4�J�a���è�ǆ ��G��}U�Or��[iv��9#��\�(2��'%� �P7v�p�!��Q<��B4��(�@�����@�h�����M�����*5�&Lé�"�T�|�V)�����������C��f������v�Id��`2�Ã�R�TNڤU�4�(�W���;Ƙk�߸�ՎqN��C�j+����?����f��\�]bO폻� v.^5E���I9��sZ��np*�]<tx�brp
9��5�+��#O��C�t_�3isζ�!z4�)b�0 �e%�V����TH��)�:`��2�����N����uI��>���K�OI�	��������pZ�fy>���	9�����[��mM�7e��=���/KD����^m�4�ߝ �j��ַ$�pzs�eO��ϱ�q�Ԉ�����jՒ�1��32I`7�"W`_�m�ky0�ez��L�����#6>Q������};ո�i��X��2��,{��y���ᬒ�D�M�#F�/'��!�r��Ӫ`4�v��y1Sӷn(�C�?��!Ei藲����������{��H�fp�����=��bKC�
<�Z����v��)>H�^`���Ј�Q�� �݄xR�y�����<ǟ�Rs♕zO_;�
�s�Q��U;��HC��	
�C��^A6QEb��HK�Ӗ34ruZ%��ORI�p��̎>��,4�C`!�:�g����K&k�[�X��i�NV��f�&��7�5,=����X�F�^��^�\Jm�#sz<W�h�D��of��{���\UOPVJ�5K�)=O��~�5��6�^C��G��U/p�����c��n���&̘J�V^��c/����z�tVwJN���x�m
X�JK�I��}��;���i��?;�?�.���;U���|!�7e�觊�'�0�[��~QCj���^S�-�Ge���?�;�d4qms[��>����)	[F�[$�ɦt�$�R��KAp��+�dy�_/Bte����ϰ��5�m�n"��[sbO��H7�l��P׸�7=�����=ÍzI(1 ���O!C����Vx����NK8��O(�|1�#�Emμ6�z��m���n(ˠ�ER�HLqL�q9.LRL�ŗ�a�p�Ѩ��ݢ��K:X�H��:l�5�F��mA��l��opr�w���X��2@@aQ3��X�̡�2��<p�d4;88]&ϗ��{V��Or��X�w�mgT��K��oɱ�Z�\y�)����x	���D�0kS�;`b�|$��J,yt���[���QI�_��h�[�u?�#^A5�_�&Y��������
�|aV�Q|�ے����H�Q{���&0%�����qN/,`���\�۔����F�y$���v~x�M+5E�h�O�)&�vA���>(+e�1z�e���j��K��] r�@���a�<MN#�������������|j%�Z~l^��4/�L�Ɯ6�
����rҕ:ea6��A�9q�ݙR2Y��h����CD�:{��� �L9tc!�|;��撿�B�,:��x$�⡊�)��� ��FQ��_�+n�Uֵ�
FՇԃ�/�
<�jN ,۠�x^Idzu����Z������p�8, $��a��ў��#�z(���Y������]g�z���^/�Tɥ�75���rֿ �YZi���:�i������bb�0ٜi�.>�!�O�=�M�$�5Л�OK/jIg�+��׿�������������E9��}���bVq�Q�P*�ْ������s1�@�)Vg�������d���Jc¿	J_9��C�B6�����4nC���0���\ƣ}��F쭘/�.�����xW�p����/B�q�ŊB���n��taރ[���Fc���>l��5Q��)�~`CD�D���D�L@���n����%,��[X�=��f�Z~(�]�#��F�gt������ڶ:s�_�+�P
l�;Z1tD�g�~T���d=�y���v7LR}_A�YDh> �ZclFǳ�C���>&rE�]�G�8���5��J�;#�S�����?��E�F]�"�J���8�� �͛���
$#�2�3�h{�A��/��U��F��	����;RLGM�����&q��q1! �R�욒@�]rA���ؚ<���0h~�2��1�}�%���n NPg�[�����>����v+�
�:0���
D��.ڳ�
MΜj'����Z�ٞ�I�ڱ`�0���le�.fbh�qm$]���Z�}���oS�cW��jJ�-�L~6NWzN��f.������6��/^u9q>�,ێ�Ta����s�'y����<ZJ����׫{j���YZ��"2��
~��C2W�����؋n�@o�����>��T����y�!M@\�=az��0�Ғl�@¼�=%F�+P�F�������!r@�P2n�ڻ_���Es^<�O`C��3�V�2�V��c{$r��g�q�e���.�P�f*,�x~��mqJ!����j�m�2�'?L����3. �>6#}o5e�Y�) �L���c��_�*I_��˚�;Y��uX��K;�6���\�!ty	�[s(��En[�Bƨx>u8��g��z͘9#��B��q�����3%Z_�E��G�xyװ��f�*����j1<�������~<X:�٤�\�hɻ盶�����lV�Jp�L��K�7�jT�+�lm��?��G�/�n8)�
'��mi<�Z���#kr�� m_��-Ȝ3�g�}ߑ�+(3�P��}"��rW\�>���p�w�X3L[�3�|c1�O�lVY���Ì5����X��l�fH�DtQ�6B&�߫�KB܆(N��`�鹋mZ6X@��pM3��%O�������9hV3��=�j��d�֯����c�f_q�^�w�f1L�kd�� h� �#[���3�/����������{��ہ!���j��y�n_-{��m���ճ���������Gk�4<���.@�'�r>Zwp���C�"/�f�M�CMq��R.��(��$�րn4��=�P�Q�1��1m�d8���i)��r)Smh
���ye�S"Gӌ��d>c��؟a��xZ� X4��l*6������v�6Js���P@��%�p�I���k\w0���vw��H4XU����jE	)�hQ:ڭW���#FB�K<`k�@\{W�V�h@T��ApB���Hϴ�-��)����?5T��M�����H���(@��᯸N��XXkK��@�emq����Q@��>&��n�e��&���	�����ږ�0{�f��q�R���)�uNh��q4XJ�a��-\+����q�<p��$UF�a��*W����E��VM�q]��+���$�l%�a|�er���ᘈ�7�[1��-��8݆Ģo��,;�E��vx%��K,��]$S�=O���[�r�1��||nW��ZZ|0� �+?����w]�bC��r���*g���
=��xޭPBy�2�m#���_���n�ʊ�H��[�'��f*pL���ä��$�p��~�d���
n�Q[���
��Dўzi�Z��%�coI����F��YZ���:�z�2�R�-:�o$5b��þA��8�O��Z/���qޟf(|�[��W������r�Uwik���*�J�>9����J�����	c'��M}�݄���rw����6͡���۬���C�:��A[-�1<;�$?ዝ��-u�3�,n����̹yЗ� Z'�@쭅�^�?	6>\��	�Ɉ,��w� ��T+��yHߑU|w�:Y���k~K�>i�"Z�:u���G�w��.z'��:9��w��Ȳ2W�9��Գ��7��h����+Ӷ�"}�m�����'��T�41�:��&ԛ%��lFhnǥFM�A����)�6')ܻ�rv�^�V�-K�:]a�&��ū׷zN)K;��`71�/�:�Q�؇+%ڛ�ā��(]� k��b4V�RAׂ��	{�Q�>�-8��)��g����6�	��Jn�*&������׶� ���%A��BN$����1�?=io���9�}��d?h���ٍ�"��6ab�/����7;�'96Be5��B2��yO����b��2K'�e/�nK�VV�ڞ�?h�F�%�y�$��	(�b6��B{��|��7��Onh�Ob��_lO|&^/D���e�}�����焸�����%��֨*ћ�ܺ��@�I��[�`� R$ov�z�ף�X���ݒ��c:j��J��2�ȝ������k��U�A���A0��A����@,x��x� �r�vr����[m'p�U��/��'��<N�_�c��׬�[�}��_�(��z:�0�w!�>�zI�7��WיQ�2+�O����ZcFۼ�s�ځ �HI�-��u8R�pAEK���4�Csܒ�X�w�ڍ�(6 ���ؽ��)���C��[�$X�����+)�i��>�� 1�^���;E�,>��M���2����:s�R¡^��0�.��[7*�|���T�(~O0�g�@I��Jm�@�� �2��_U���4u�8����>_5$p4��t�rPc���t�VF�קeL=����u���6������ν��+�߹�Oy?�i�W�����ۅ9�B���V��Y�{|�W�k�G�D�P�7ޒ����~�Sj����&OC|fc_}̱�_Q�0��(�;��d[�9���Oʱ���$���=�[bi:ݸsn�l�*2�<E}�?'QXE(��V_�N]�C����؍�G\���Wq;C�屓>��Nr� VJf�k:ٯ<���R��x؄�M���i���]����q�v����B:�o��0�u��:f��E�@���v$���]���+�-Ls���ڗ�/���}�&�b�9�`�K�2R���+vw�US3+��������O�Y��YP;@�}�v��/�(@����-�^> ʒ�? s�l�������9�Q�ץ4�7� I���|�鹱�|b$۟l4t�Ih�|�O���f���7d�:7��љo�á��_�r<pN�m�����@��ݣŧ��$��u'I1Z�@�e��U��n��C��3ӥ��ײ� ]����K�_,}�����X��Z-�a����w	�yy�����_�cQڔ�6�3��������\�a�E�F�:��o�����/�+��u�䂤Rs�+�4�x1�V��c���K-��B��#cUW�$3W� z ���M�RP���C��ʏ���J���*��-hq�ć�l0w~���`q䃜{6ԯ�q{N]�>\�=Nd�Hx��y3���T'j�a�@bH4�?��E�h�El���cX�<�H��ƻ�)�ŵ�k:�M���_��*Ѷ\�Ws]h��:#,�x+ڕ����{�}���Q:��.oZ����׎@O/=h4�&�LM�z�= g���3z������+ҹ[	�:�|p=K��ó=0Z�q_<|Sl�/ �I��ϥҍ��s�5�c?�*߬��{1��g�0� �%Ce�uTe!_o�Ġ���k��x�_���a�Ѩȅ��Ӗ�P��b�B#�m2X��{�Yk��N]��&Q���+�
r>I��+�5}6H��J䰶ѕ��\��Z&��� �����`Z��܉�k���g�Ͷ�7ލ���!=��ڗV^+�>����~9�Djש�q#п�k�B��T��J��C
A7u�|-�#g���l�,�>���YtIyb !���$��t1z����.�+^��`��r"�2�d�,ez��-=�`O�P�_��9�ǣeQ�(g�Y��W�	������c��pL��#t��;.R��X�����O�F5����E}R�D�
2%x���
G��n]���|��Ll7`)B$tk�p ���-͋L{mf��u��F�p D ���w
xy�����ƙD�H�LGE��yx�s�[מ���K��	 v�v�,t�u���FoՍ�ˊjy�1�E�(���PO��sP��+�Gr-݀��2�кvy����\^y�u�gLH���"���H�d�$���-@?�"f�e�_J"w������B�&�غ�]cfs\��me'�z��R��� boW邟��|�����~�Ks�f4ؒ��T*�h;d�y�$@���*S�t�R��6yk�a<�w{gRȀ�'I�k��(M�|�O�2(��[�F̆H��?����<$<��&�h��aRbW����=�#���2����@/
WY�2��uS �F�ǿ�՟RWG���,�4�8$�beO`�s��Ay�@�p�dQ��s�VX�E�4�� 	n v�)��\&�!O9^�λf+P�I\�����gN�選��=B��J#F�*����Z��!F�\n$"��O �	Ӽ��8 ���F��!Y��oך���Kİm���w-�_�"ag�����~��eb���ۄ��B��9.6�XN�����ˉ�0�4o��]�b�4.)���á��Ȃd�dA&�ǉ����H�=�BM3y�\y��'x�B�Jl�Ýu��d˶��l�+*�x��T���� юD����h2�P�t��Ȱ>�/���Y갭��
gvH;S���/sc�ki5kkI{�-�] �>�5��I�xw���ĩ䇤9!��RoHJ;����>���7E��:���}��ꪶw=��&�\@O	 8�-�ۖ1F�a�`맍{}��v8kv�p�C�8�[���Ӕ)�Y�ZL��>��g����J}�7�5���z¥T%W(3�����y�^�Hc�.�s)�ǹ+�mac)Ll��%Q/'����S
���m~�[셾qm�g���n��OA, ւ�\����-'�uH>�I3Yu����~�ֲ�_��@Z؇�*�:�&�?�3�-��1�,����|A��!Kþ)��\t���Ȃh��0��t�?EU�5�$�HK����Y`����DSzgKf�	N��̟	�|�4��K��+#� �J��l�7��3�sU{\2=ٝ��UCOTJ*��!��0M�BK�/���X9�+'J�q����d��f��7`�-F~�\�|����]*��қ��ĩ��V�
W<�hwѼ�.���������h�������-��y�&�_�q�(t��x���h�?[T�7�cC�y��<��|��d��1Ӂݥ��B�`�ď�F5E�}���C�ͧ)�$�%�h�s�n�ɧ@sч;��"�e�A�M�;���^AE�8�1��}���¡�W���^������U�����E��%��`�k��Z?�q��(	����y}��|=���lT4�I�J��`��U���Sx��l)雹�x���������k�vE]!M��~(4�Y�:|pA��"_��6?2��f�w�����<4̓R�����Ɵ?u�͝˥�����!���[��V�7���(������v�ViD�@�N�4���-m@���3+`���͋�������l �q�pQҌ+(#��O4��U���{�7Q������Ÿ�o&��Q�Ǥ�t���Ekz�KCh@���*[li����u���3�kI�EsY!9|��+���4J��J���o~�N�t�U��X}�CVEvp��	/�^�p��H33�3;	�O�hZX��x0;"��n��a�r�n?�9�s�;	oۮs�@K5[��3W�"�$~Ĵ�g�a��Z�j:�W�u]��	��A�%,W&�^�>���W��Z�Z�-'rF �Ԙ�&��� SkI5��~8D��7�� �����wf�X:��
l�q�$���Ċ�B�ǋ�|�Y&9J˲JJ;��	��%>��˶T$<�M�Rx�WS<�8EHcu�}���L�2�-&r�U�hk� �8]��M�N
��%t��!ٝ�x k8�D��4MX�8�V���EQ�z��(�^gu�����y_ �F�����|<X�A
>/d�<{��i-+t���l�g�\kiWV�C���]��7��7���
�C����G������a�9\Ju.1'8��^��[�7圱�"���{似F[ĝ��+�W'4�]����<S�����W-Jay���U��Py0�(D�/�K	{����8#��Q�k�Q�mԈG�HD�iἪ�M|mٞ/~+��+s����ՖjX�a��T/w|�����2��yݕ/".�l�B�H�Rp�����ʚW�������A��A�D'��KT�yx`��ĥb����vQo�{j6�x�dN�P��`�e__ݾ0�Gn06��Q��9�d�Pg�3"�r1*U��MY�B�[jQ����%���m��~��ޜ�|�m0v_�Hj����m��4�1	���8�bQ�W��I��׸\�M�'�?���b��tcC`�]�hz��u��Zޕ^�:ӆ�tI�f'��3��.@�������!="���!�ʣ�]J��`�r佒�<m��Q��h�7�:c͒
�a�"~���Y]��g���!C���Y�V<T���v.���j���i�����<[%�_>d�m��T}���A9���j�h�؊!�(n�	1�D����"A-k��ȑ�.j��v��3/[��d�v%r��/иW�f0����.�ҟR��n�m��9|�3���N^���e���*c��/�OL?��I��un8�ꉽ}Z��X�o�����n�9��®�&�	�g�[#�k)��~�=�i�
7�(�A50Әfx��V��r���n��`�_"�zO~�K�����ڻԪuP��{�a�(�����k�������%_�rԩ�YE���A��C���-���BOGfd�˒�f�Ն(��xJf
S���ZY�����Qz/R2���N�����Q�`,�Q@�-TV�Ht-��J>ؼ�GRs����i9}D]EӬw�G>�Ɯ���x���w&I��x��1��vʺ��w�D��$s�����2k[�9ۼ܈ҍTKԷ��ק�{��ǽ�6M!>E^��mdP��e�n�<SYI_��NM��`�(Z��U���\�(�l�ח����T��p���̔{&B��=S~|��
�y����Nqr5v�z6�-v�_����!�z�O�_�|G���;|�=&����(�B %k;�:�����T�d���ؗ�Hn���O�H�^��~�j����7�;��*f~h�-��{����11� �Ѣ,���N4�٤2b��S}􋞐��?�4PW]�0�?Wo��FA"�lC�6ӷ��&w)��C=G�(^�|Na{x�M�s^���B�b��7��$`��sC��9�z��0t�����X��mѶ���Z�v+��#�bT�'s�`��w>��(��y|�샐�sJ �v�r_�j�o�/�M���G�ہ-�~%�7��!�t�hzRX�Z�9E&|��ɢ����v���t'Z+�}+��7�p�;i�u�{��`*��σ��)��c�I�<���p�3��@-8���3Sr[ܢᒜh�s���<�B(��V���	7zj�~�7"�K��Ӓ�V��љcr�u��Z�'�
Zֻj^����q����	�nȄ{sY��OL@��]N��p��zL��t§�����o�t�@�a��Y�˻��
L<m���s	�5E��z�;�����3��{�~1��ko��`n�/�f�	�ի�c�\�p�=�f�^R�V�$��]5���n2q�|}��S��$�j!�f�0�)ij�X�8c�d�>^�l*�I�K0�Xv�wόo_h@-
�%GB���qA���r�)��;y�W8��b<��哨L����QHX���#G�?u��8%����	�!P�r�`���~�����B��B�dH*D��\*�� ��2Fn��R�x��ٵoj|ˬ"��c+x�ht����-_��G������C0-�K�D��
S�D�uc��S�%3�壦~�!H�5��xH�:	���X+u����9� J����@ڄ>Q����s��ĴolwB��f���������� �Y�"��i_\�L^h���b	��A�\�^8H�a�o)�D�f�|����]T�ɳMV^Έ͇J��eƇj?��c�\*U?� �ǹۘY��GڲV ��H��^"}]�KEK���{���ȶsW:ga����;�묏�/�)����`K��w$`��Y���=��XPӉ��d��5.�O1$�{��?��s�"U�G?O�B�6�����W��v��;�p:9mi�yP�o��'v�a�Q�چ�bްB�mYTu�1�@�i�Yh��g���!V��M�H뼉�@"Ը7��<ju�:��T�m�=�fB,����3N���g�|x{le���瞾EB�d����4&��bz:b�z�p9�)�'��zq*z���~��J\bߑP����z�	}�G,2�j�|�����s ����Z�H,�Ny�a���~�:��a)Y�1������4t���`�6��3\����/d����x������s��������a��"�E�]�TL8�Vj��K~ h�\SE�P�(���^�V��0U���Yz+0�/�N�/\�(g�Rm���[�mO���7�,^�By�I՚��YF�i��B$�"lhۤDp=e��|uX���KcJ P�ܸ�0~8iu�n� @c����J�$	��Ϥ�����J8�_���T<[{5���[�(��_υOZ�N�s[x�]Ln�p�OVVph�V��Nd#2�_��S�-@%�z�2 
Iv�Ţ�����-��)��:	��}꾥7߆�Y�+Y	о�Th�����ܢ+����U�����
8���M�b�_+2
�#��+���WYx<�ód0�^�/%�|��54�If9�4!L�X�q._kC��>��
���� RJ��[�K�Mn��
�Tj	A�\!߽�ۺ{�]���ȏ<k�Uڂ�N<��<4�D#�����M��ן����ƽE�*3}˰
HC�H�(�2�����d4��1�EoS'I��J��|��I{(�z1~bI����u!���D���x]�s��JA��\��]}:\�c��A�LR�a%��&kb��+!���#���>UWƋX�Q�.&��D(D��s�pzV:�<�f�t�E9n���<��G"�ǃC�U�����ѹs��f8t˅W�']*���;�EBm&�s�QV.���L��`0b^ڝb��D؁9��P��LH��aD*�:�$2�fԋN��؇�C\M��T�ּ����O����v��W�(��i�X��:�\��K��i���Ri�o$�8�>������b��+`F,}X��1&�b�����&&R��>����FA���7o���0�G�����r7֚�G<͋	�ҏm�$��o۠�ݭ>n ��<�xz�����/_�9�ə��9ƛ�Y򗬗׹��v}Z���olX�����2f54�Ė��r���6
�b#,�2���]~����������X�˖@4mJ�#��֙�
��kC�"��H�[Ey`1{�F�#gPTބ%�
�ޔ<��7�-ݷ�'�JѴw~e�\R����ї��-�列���R) +�/٩�	&NB����&zk1��)�E�zJ�2=	��[	��/����#<�0��\��sY��ӭ��J���z��XG7[O�,?�3���|>�=|���1��9�Δo�X��9]a_���?�ݮ�c��ZA~ю�P^s�y9r+sɤ\=s@���ԨKu�H�u�k��!�F���7���V=�`Q93|68�~��7����ǳܟ�����9f�}̝�;t��Mx�NԂ C�9��^�f���{>�X��WRA��ؼ��s���,�7��[���	^���⻢�D��^�ڈO��677�o�?=�A� KJQ6���]*#;a����D2�:�V9�[T�<]M������>f��u>D���E�n�R�?��]���LNw*�2�%�࡬���>��R39���Y�|��\����m 	Ps���|�.CB�l]�B�a]�P��<�p�Bj,�r�r������l���ӄӔ�D!y}@�Ea3`�/�r�@i�����w�2C��h����S�fՉ@te�w�疟�?�O2�}-F�/�;�]�ϻ���F�Dzo׉�ר3Hl��C��<���2��^��w�x�b#����N���
x�9��Z�l�b;<��-%F�0�{�85E_e3�}>�j����W�6�Z���"�I��E>�  ���y{�˔��˖��h�7&�A�5�O ��z+bEj;�LnV�����V�g��x�+�˖��}mw?\�b�x�A�YhV��yI���X,���b1�^0��r�$Y	���Q|�&�KL'~�Ve�[˝4�Xl�=[˞�UÝ��2�K(O���ϣ$d�E�r!haRAE���5Bf��d�G1`�z��y�{�r�bl^;��-Q�jyפ�Z6�wz�/����^�FX��Ea�b����.���Y�*׻�cچ�+�كr��EH?��~o#�+Qؔ\��KW�.��5�-$�5�]0��7������)ඩˁY�X�����"�l׾���A��S��K��	/Q�1�#/�������yj����dӷ�L�����|����|��npą>�#�����/f��{�su�%�ђ���CVٯ5��4�4h~�
Ug�B�ӛ�Y����f|:�jB��ɷ4��="�"�Y��G�>�D�Krj�ʿ�G��[�脭b�#u+B�>�C��l��I��@�O�H�bx�n`��	3x����3F��K�^��1V&p��N����x,d�d�}N���-cV&g*@R� k��B�|�jq/ڼ~hGF��J^XqI���mre�p�g� ܱP��E����br6�!E�\9��֑�B�d���y4�|K�%��L��C��H=N��)�(�����\wg���ձY4�>��*K�3��pm#�������ݖ����L��.�g.�A*�P���*+��B҇�W��K��)�M���<nX
i0C���w��^X���g��]��X�����O��/� �t��9M�[{類y���/������=:�)����ޭ�%̴h3���\�슕l�~��� V��oO���F���C��q��)H'�DN����F�xZ44x�*�j�����`�^�b���W��FMN>h��MM��dJ��6�2f�X��5�E��
���8NxQ�����
�F�c[t[5����E0�ш�y�Ɖ��[부�Z�7	2;B�>�C7��P;x1����M��z���	s,������3��96M�ѧ��rU�p!��lj�����Fk02����A��;x���W���З�`NpqM�I�dE��*�[�'�5	�	1�dQ%�w�!sZ�xXƍ�7�?�޼��81���Q�H��,�����n�W(�|�c� B�5��-P�|�0X����_hn��l��B�Yx;��<�`��DhgLR�i�z��9�ms	?B3����e�cI��o|�%�S��?i���P�6�X3�J4=��0��r��?*�AJ��a4z�bv㱹���yo	\��D���G2U��2��G����7q��d FN�1�V~{$nX�<<[�$��S���n�R�ѡ�m�[O�����t�Ҳb��ˤO�Xt��!�FW�QR��߰�M��!�� ;��L2�=�~^�.�yc�2}�������(~��*E�t�-xt�;|[_K��->Z[�RY&(=�yv�Z[u�t8����C�_���3jy�������uP�,K�k9�P~o���wI!��њ� 1�J��{�_�d�
�b��æ3.~�7�!���|��x+�����m��N��n�'W�×��j�dto��.�)�`��Q��#"����"x+�I0�c�C�U����������t�c7�Wz@'��  ���ӿh���T�H���Dl����7����U�Ĉ\%	�3\\�ͭ��f;�%�v`7f�x̀�M�F��V��xp��Ƃgx����#7�0^4���K��tKR���sBU�&v�漁2�ĺܺ��2_Xk��Vj� �\
(�t��t��*����2uI�8��Z'\�j��45�dD��)�$��XD��Ü'�rާ�z���ȶ�B�}j�P�k��X�9��R/ɍ��<8���c�9[qD�\Uۡl������*kӆ�N�vi���¤>B.����"�`��p���r%�J̿YԞ�p�rd�+k:�5N�
v�]r��#4���z�s�@��9�\f���^������O����B�dЫ:%��'	a������	�|X�>�B�9�m���7��fe���tÅ ����7���%���Ji��c���F�Wge#��ҋz��t,O�����
0
o�W��)-�02�v*Gwycy}&�#����7���l��
�7�pj0�_�r�zF�x�E�=�=h0�l���C�4�q�5	/9�W����P3W�	'��]4��Q�V�!&�~��:!SG��=�b;g{@5d������� ���h���'��'1
�9ls1d���k�3Y��_�f��`o���"���i�z@���RA"�;D���(��}��~l���Z��6RUupX3je��B�B�Y�k�����-q�Ii�>i�l5B�X����s#Wfܖ��
�^&i��lc�ny����-7��e����;1����a�%��/���S�>w�&T�H��K%]]���'��¥�<���3C�ո�'�f�M$�HކUt��K�e�wy8�L�h��w$M?�����t�yn���A-x�I� j���9�1HbP���]���hT"�)�P��-��g�m�x���]��a�Mq%P�H�p��6��!-����c�Å\�=�O�����r_9�j���G5�cq��i�	�J��aa����- R1]�$b��EX���{G�Q��mc,bϓNv�D&RT~_*�sj�Kp��m6k��PZl�Un�Z4��	�]��y��-Bw��x�RHL��<��sB�
o�_'6y0D�ID>)�}��P�Ô@���*0�co�x��eץ8uiU�w%][�7�і��!NK"�Y�����+�r���l��Z�����o>ݐ����Y�$6�s@�s=|'�Ŵ��_T8���F�2�Cm�����=ᡶ[_�r��>-�f�j�����
�3�?�ɟ?�j<�3X#;�&{��tP���m���Q%^Ċ�d��[e�e�d��s��i7}G�� ��v;��� ˂�ys��j�)��J��-ꬱ{���hN���mF�/��\�BH	{�voić��1��	\P�|n8�(@��К�S{�>MY��Y
fƝΨ���&-$pFf����s[�M���ߜȕ����]�� ������,6L���D��!~ۘ�Re]�>@��'˴��J=̐~a��`��ށR���A#�.�lKר,9����>E��mB�ų�g��l�1Pl���n�,37�s2%��|�=�Ci�@.���7bK�q8k�����W�E��r��x)A���걫d����|�Λ��Ոؿ���C�޶�6e��I�j
�T<��X�RN�U.�H�o#
�L'��qoQ�Zd|fP���:=\!�X���s�����"��J\��ø��q"O�A�rps)m9�f%��D���|�D�>�	B�Iy�:|g*M�=�d�$�G�J�~ns��?�Ft��N�7~ЙB��2�󲅏P���OfcRw7>�Y[/C�4x�C�\�Ч@+�!c����@O?L��$���j%5���*=^n�=��(��Y��HK4呃X�*MU8��X�*Xs���0��,��a��֜m �ی ��h
��ު�bvv�������v�Vg�#E���u�!����s.V�/��J'f��y�$�9�����7c X��^4��"Q2:G@�����	�?���r�Z*��іh�@�zV�u����p�b}�aQs�
-�EuQ�#h;Ʒ`/�#'&�7�� ���O�Ѳ��7gxt25�.�I�_U�-���6W�4�^OJ��Փ
�+��������1��NJ������x]
���&Đ���*�M�oRS���� �.�E�h���t�M��ot���R)4�K��l]������%�1��V� C=}��lV=���fܵŗB�v.u���k|�Ѹ:|Q�Zٔ
g�x)�\�3�E��Oʘ1����O!
���m=k(E$7x���V��T+�Pk1F���Y�b��*�B�{�[?�J�	��������:��.*$Hy+H]Xt�b�E:q!�T�5���m-��am�y}�u�S�����jlӮ1$C&�?L?�z�Hmа��r�1�2Y���w�����n�\y�x�����/�����~��>U��o�����na�t|�٦|h���� ��!h�s_e�=z����%��������/C��O�;��
�Y��l{���'7�N������1��Ӂ����~l\��,�e�p�~b`�zu��2-�\�_��2K\���Lg�p��n�^~��!�
 6�ћ#���>B��cG��1y��$��G�P�nPT��&C�}F��{����Z���機hP�$X�վH�/}������_M��c��݉8U��i� ���1�3y�8g��.a�O���	������i0.��ʟ��Ho�0���
�
����k�ȕ`�-���+�P�bc����HP���y͙�w�bR\ƍ�s�;���=اk�pr���C����(Gܧ�-�������s��%*��"���L��s}���1���N�W���l����J�J�=Ú�/9}v5�"A�����м+�DN�/F����0� �v$`��&�:��I�KC���� �9�E�]KK/�y���|j��fb^��xz�m��0ݶ�*|xK�6�0�W
���@y���E��mV[�A�>�f�a�>�:�0�"Ώ��S�c��F�Č�w������J�T�򣂗���͢�`yo�P�⎰ ��'�W0�2&��`�Ή�7��[��l+g~V2(v��F�6�;Q�蹀̑bg*��@ܴgf㠪QЬ�r��H�2
��d �ćߠSEJ��1W}:1��`�D���Ww�
@�u�Fu��Ѹ���q��S�f��"U�����o.�1t�}@}�[S�V��+�6�X�\տlik��
\�s��ABP4_�3�so&��:2y�=��_���"�/�\�$�j�6qTهZJ��1�7�
�ԛS���Y ����}3�Q��-�uU)՜$���Y��*�>jt�H�K[���5^Wn�N�~zA��`JF�=��_�❛�)ܪo�i����&�L{��!|J�Z�S7Y4���{y��u�:}D�sJ׻�`�g��.�̧g��6�D�~�UfSrk_2pe�JT�yb1�:����*뉍G������E9�`~7�j�����)�<ŭ~U��og��gXOF/āK�t��in����+A$Y
��a��S�B` .W�� �~.����ϓ��^!7m���5� �lk�ѳ:�ٰ���X�9��
@ŀ��﷐y�ף㗀H����m#
�����+��W�F��|H��A?:����ߍ�NCHh'�N֞�e��}��$�W���C�Y3���Ҷ�q����)	�&(�F�جw�������,0���Z�!{쯽�$�im��k�c�W噮w^R��{�̗���}$g�sj�qt����%Jb�\��I�wÎ���G����n?�!%���@tJ��%j�(�����[�_���g��-��[:�lI����56��~�I/�I=Ҽ�i�.���P�Wot�KG����L�T�2^W�Z��� _�̑�F~=�?�Dp��\�*��3�k����ҝQS	S�X�ͬ�[	7PIP����?/���Q�Ի�k�i2��|mȂ@�F:�F�ל��#�]A 志Q�o��MGM�"�''��b����.0��1*�J�oG�B�U���5�y*|��K�yΡo�uh�U�`=�L���PDE,吥E��	�B+�S�c�X��ՍV:Z5�t��u��������Yq����2���P�� ��i]k���,;yqM�֓$�|�˶����K�z\�����dk� �n�]*+]�)'W�՘��Th~Y����K�ObeF���-v�G^��(����qe�d��#�8ۡ�1�v������𖛩�ݛR(�B��Ή3��8���ndt�^�y3(R|"YH�z5s��pE���)��yeƻxe@�0م)^=�yY��m�tt>*R�cvx�;���SC�a��

�>p��_�5�q��)?����;�b*�%��cl��I^	E�/�HC����Gv(���Ӊ��s���'N� f�:��c�o˷���^:4w'('��e�U�K�s�0�8�u��|�V�W,>I1��9|����J
|�����G8�d�S�˞ߘ��٩�AL��q7� `-� yR� ��a�p���@ңL�) �Ӝ�~K�
�?e��?���%�Mf���Ucg�b�������w�U���rb�_��{�e	��h�_����Nc��iδ-��(����_��C�����7����	>�փa��mi_�h��~�C�Op��zz5\��Ϋ��T���,�j��1 ��r�����"�ZT�j�/���b�y�{RQ�!�	-CPF����������H�O Z�[��u����-�`%[�ّ�e{� |��q�S�&����2o
{��L_�}(����"���_�Wt4F,n�*V��2	]Gu��@X�vX~Wբ�WW���ą0�RA{�~Ȍ�]|�rEJt%)h
�f����U��xf�t'����uKZ: �����"�b�_��@
 FTJ�RF�p}(y�=��e�t��	_a85t�^������(�up䄎�sx��Œ��zԲ�;�c�����gǋ��ʩ���Nd���.(W�Rk���t��x^:�V!��9'E�nz�`�;c�xN��;g��Cs����F*m������~�4~��;p�^[ِ��(}q�rz{�j�@��6EI�h��.���T�CT��c�z�@ શKWz�V�̕U�G�����^b_B��a�>!�L�-��BIQ�nB�h��&�D/Xi���dH�A���5����d+ �-ƨ�8�}rJ�o�Pև��>��6��#��T'���|{喯�7�빳����ڡ�qdky�q �@�pL%�p��@x����CO�z�VJ���N㱟�\���!c��>]�_��I�_4l ?���^r$T��U��΢,.wz����{	�K��6�AΘI4��f��i�t��O�׆B����hя�W��m�7�c�D�'�ǿyV~��ms	M�+nb�k�@�1b�_d!+�Ye÷�a>�p���Kǚ�(�q�S�����q��7>�n`�m1xR�xƚFT[$��)�����J;����UPݞD��_�6T/���9��O1 ݡy��U��ݘ��2�{���_����e�7ķ�����z�M3P��HfSA�:��\��_C�w?����r.X=���|����ѩ�����V�>���7�^t���?�{#���Z��	�BʪC�d���$�P����mW�ZuHx��`��~!_������ѣ�)u��N��}�:N���u�!�*�,;�ZZ��]�F�/KVɚms¼J��[�Gl��+�/e�1$��������U|D��C�%��a��(:��vH_,��λG�m��nf�,S+��d��^b`��ؑQ��x �}�-W@r��s I
����qe�qҦ��"'䝩^���	��6ܭ�Ѕ����w��J�_�n	�b�FuC�-Q�µo�D������<��3Ь���: 7���"�d���m�Dy��J���]f�&Z
��-������Lvo���90G�Nÿ��]Mb�1�%!�c��Bn�W�j�r5��������]�U�Q'�p��(� �K����7*Ԋ�]~Q����4�+(qϭ��zz��H����a�m���#�u���n��v�"L���E־��-��=�3m_(9V���R�l���'��]P��/�"���v�0��Ζ��.���5�������AđZڸ�VB�6��dA�a ���pT�J�!�m�t��;ĉ解��v���� ����]���DQ�8�p#K��F������'���͌;���2�}��e�:&W�~u�V&ze=+&#y��_�>rgHk?��ǀ��W:�"��j�B�Fw!���3�E��Қ���*h�"5
0~W�&� +(�n�>kjD=8��5h������龲��z-
�+��K�{��I8S���&���̺/?P��#۰ԼU��+FD�
�
���;���P��΍|^�{*Z�>ޅ��_�}l>�[�uE}u�S����0{�qiS�Xc�{��+�|is�I^��G]D_��7����)r�S��(���aE��� ��kp�e�g�Ǳ0�Kا��*S�L���2ɀxNo����yS@6	8��|ɤb���d\�f��2��4�{,�x}�ks*\�OIn|��H�lk.��:�Ƈ0B�� �E�l��Tk��Y��Q�r�ם� qSc�	��|�����v�_՛�q�e��HeP���1�jPhp����P��#a5����P��86ce����"q�q�WJ�&�I b�-�X�,�z��N�6S3�ª$��P���$o,�۔_[��������;H�����,��a�0ńuh���ɹ6�^R-���yCQO9�SۃK\�`�d��i�14Y�{tF�ҹ����^�����;$�Ba�"�A�nUT�J��t˃��)IGa���������K1�P�ߓ����uY�3K��f�Y<�1W����k~�%�\�.��L�-���D4@	�¿�am�&��8�`�8h'��S�����fmf���Țs���c��e[�p�H����N��_j;�D��w��ED�A#�́�`wu��0����ͱp�@��%>酔YE6�?u%�j��KXx����%n{�.ji�.���>/��Q�����<s�{y�!Xk}T��c�1�@�)�&?��y{����w �+} �{ ʭ@�n���=*Ċ��̲����,\i/nę������k�J�BE�r%��#��@w��.���}�@{DMT���?�;j��NUL�ms������x�J�MR�j���_q0-:!��s���j���a:Ɍ�pnj:�m�0�Rb�}eW�&�]�i ��J��� ͞D�"���	d�YR�������o
F����ٷ�j�E�<��D���x��x�S������_X�'��GR���U�΁|{=p� ����[���ɯe��z�y���T"�3.���g�����w>�ļ����)jZ^V�OK�#Y>�%L�%�]��;_�b�dW&�̶�>B��qw���!\�4�vt�9�zj����*�kb�b�҉B��
�������bY\H������:��O��F ����5[��-؃���*is��_ޓ����as`��:�56���4�+y�����ܵ��Ʊ�T�x�1�sj��h�IۨY�5��li��[u&Dw]�(� �P:Ǻ�\�=|Md��yә" ��a�.#ǥ/S=�Jq�����1����b��|��dr��k����I���]�*n�;&���AJC���\0I�����f�CVhz�iBC�Y(!p�P�FjZX�U��<��JpO�0��x��yi��y�b6��� C������N�N����- sϽSxB,�,UY8ü�g��9.������"�ň���2�����6�,q�[�5@n�$o�^d{�z�9m�h[B�=`�1��?rX���� ;^2'#]��C�	��˙�ni�nlJX��xsԖ��P�ɒ�=�|���d���!gڗ�YAJ�o�P����05+	T�7�@�i��M�kR�SYhˉ��jt	�;;�m o�p|�C1v��r�Q6&��=\�6.��!�0ށ��6B9�%mػCb�E�u�G�T��7��L�fjo�jeϦ�Slrh��n�n��_�A2m��7D�	
�!k��fJ+��r���2i�.`�t�o�	1�?�B�@j�Q��U)=k hؗX�#�[��̔�8�m���	@�9D]��7�@��H����(,����aކ��}�{'1�{p@&�8_�eQ�o�rGB�փ/6�ߐ�B��j�S�C��q>���|9�!�(v�3Ȥ�t������Zq�/l.��1�#b�v���gj"��Q���9���4��P��pMi�abx)��Ш8��{J�WN�q�S1)�F���/�㷳�(,d}���}F ��F��E�Y�M�$t%Y��P���A�RVO0Rxɀf�Z��he/(��~�l�o흷�;�=h�>���e�S�nJiŦ�v�{H�7/�&-���>���qW�wu����z��O0M��{F�h��� �Z��Rv/hֆ_�l���?r�^�jF��yk|�81Q�C��6X��h$����
ɬD !�e�<P4*T��©FbSr�|�Z_
�iE�#@���8@,�<�K�Q��C �[s;��!����n�ؒ�}�3����N����{��G�=r�G��e�؛wa��+�g��C�W�q�'A�L��]}�� /*z�vao�+Ts��RW�Aw),$X�(jӣ(`�G[����W�~�L���)����,ޞ��i)�*�����U��{L�hqaKWV��Mf�Kn�Ã�9j�q��\]3��^pg�_����&��tgg��}�� Az��?��d`�C���u�B�5x6��x��
�-����tL)��"<8!Fۤw�!{��˔7I-�*�_�5Dχ����`}%k0��h�^s2�,�<����;z7�`�|]�q	/����Zvob�Mm*c^YZ}Ub�vt�V��y�Gmw�-�~W�+>���WӜ
��	(���ҭj^uD���@L�뭓�;�������f\ ��o3�e���]d��bi$
��'޷���%�c撿��0zǉdͅd�/��0�\���V��P?H_$w���+��t��b�V��N�*)�xڦ�a��S�\��_<š=);�ш@���N�q��o&}�i4zO�z�1)��(��������J���J�tU�-���0�>��f���-=�&h��*�����z�DC[�E_�q�{�������IA�x(�T+l�zx����ě4��2x�JS<�2"����mX-r*��C�Bi��<�����4�]��<sF&\�d@SHJ+�� ��.;���2k;��_/�'4�@�H���]���P�?��Zb��`��(���׶����x ��Lm��7h�o���ߏnԼ� ��Q�e�F��.��";d/f�,ͮI��\�܉L�}(��<�S~\�VA�`Q�q����c���n�y��k�01���"��e��	4�>�T����,ceގuvR��wo�j(@�Tf��:LM)1s#���|�ᘒ�і��2���L �����Y+��e�ʤ_N��O�8��6+���5g�Pz�� ;mb�m����Լo��·b��tɵʓ�:��ٌ�#�*�x�P2%|��Y��,�>"����ja��:xRy���T&x3��➽T�gp�%Ui��H�,���풆��l�ַG��BO�)�H�Ypq턨Ӻ�	��"��&���V#��}G��N�e��փ|ɽd�����=��(d}	o�ڭ��V-4D��:~�v�L�i�����w_�x�,$�L1�PU�w{&��Aɴ)l�=%�=�};x<��耄88�<�s����zV�����5�����_��l��c�u h?'�/q�ډa� �)K]P��j@�0z��ml@ i�1�3�R��(�I�U&Ʉ&"��F�5O�A�8����� ��
/����<�G�j�-9|��9z��g��viJk�63T�揖�nN����	��"�z�7���H*9�N<�D�21���#&lA�^an�@����o�����g�L1��>�mzs��0���(8G��[�=(<���P0G}H��V�L�l������]Z���M� r��x�aA�J��C͜>'6\������RӴ.���=cW�̼`m��D{�!4k-:�j�1a��MB��[N����I?�����r��c%v�ڌ���_1�����_:�n y��M��5E�";�6�c��m��PNH��--���$��%��f�$[� ߔ�����������t���%;[�U��'�9�`r���k�=������!0�ى0 �+�C��V��~"+��<�3��@k�0�� 6�\ȅ�~:�}��7z"�s��� Z~���Pŕ4F�ҵf�.1S#E��, ������}�9;�ݖp�~z㡘P�yT��o$�q��Z��9
�Ԋ��;$�p�=`�ɯ`�?�#|d�>m!��s��,���.�ju5��9�_�~s�俊�N��\I��)*�њ���Q�d�����A��x��W�]+�>�>/lē��a8s*�G�+,�+��h��g���jk��vj�:����ZSO�3{ʊx���Mm�(��Љv�����1�����#�fhޘ��4)T�� 9��Q))o����!Au|Q�`wH�%��17A�{ː�dƇEc�H"D�ᖄݏZT���r��ص��yr��nM�I�m�U�|YGf�2��pBp����xd��S�Jm̚WiZ1$ܜ0�7��M �)@ ��?�{6��_t�f����(��~�L�qp67�I%0��s7� ����⩎9H��ᥱCx�#�����c:��X��rW�`���tl4
:[�ɜ�HSh6r�2�?�T�����<��J��h}Om.uQ��n��H��y	�̋f�≪/�@C�$�UE�D�A��\`rr��X'��ZT��C��V-@���lW��ی^!R���N�eM�[�>�CjM��r�
k��؅�uK@�����K/��K<��ja����Aa�t��k@^D� j�hdշ�&ou�8C7����*i
ҋ��"<ٱ����i��U4�|�9�S�fMu���$"�N�s���`2�9�(�^���g��Jޓ*�����}�z��1?�*�C)GX�IhP�~x&w������]�tn�@!��d�>n��E0s�VS=��H�T6��� �pA�j�7��DG@�N�}�EH�1_j�lp�50j�o�i"��8������QRF��x�Z� ��s�K��~7(�Q��@��Wk}ƘU���e{���t���ƞ�k�:�	�qR�tћW���y���玏��z�1�'#�b]~7�J~��z fv6)��.�k��f�!�f�k)��W�Lb}������3��Y��ǩ}?z"����
����!NR"�~�&]u�	;y��PЮ��Rkv���y�~>c��l��<�P�FA
�i�D�чM�h.v��R���8�i ��m��|�L���i��:o�{�ů$��vmX�y�Z�lt��~_����Y�G�(\n
�n�:i9)~툳,e_�ݟ$q[P�v�u�y4V�M��mL�y�u%3}/I#�s�`�{�_3ү��;�@���D�6o�����k"��q8�?�Ɛ�R����P#7�y�͠f{�8��U���e?��#e�oC���>"s�S��WxWY�ރB ˦� h2�NA�ϝ���+!Ä�R�����`�[��'{��
י��io�m��S>F�n����u>���qԠ;���*7%|R��;l#��k���3HA%]WN��O�!� 3&���.:iN��)UB�YG �J9-��1��B�����:����pCX����P�3j,��{	!1(�~4����:P��ݽ�v�S�����'�����'p �d����J��[:���И�8�Wd�`D"\<P��XR����qP�AÚaZb���J�D}s���k9ɱÒ?��`l7bZr�n~ѳcӑ����H�p�v�v,r
�-�7��~}�thFɋ�$>�B�(�\?;m�@l	=Z�mY�&��!�,%و�0���)Xs�Q� �wt��_�Ҡw �e�*`�4ҘV�1�e"��$���<Ү2��v�U�P��k����X�kB�����H3�6YT�!(��������9Ic3�&觮-�nР'G��ǐ�%�p�v��"n�VO�c,t�κ��Ƒg��<D!�_�H�p��M�1�1c�5�/,�O+_�l밸/���S܉�ׁ�Z緓�ԃ�P���]h�� $�+z��s�:\��s+��o�Nb�Cj�ޗʜ����)���CblK��~�;\��#�<ˤ��o� �e�����[6�x���<���e~�ؕ�]2�� kלҠʾW�>�37Q j���Ӛ���j=�5��X���TR1���KL�z76A�>/�.ci��$�t�~�Tgb����ztuj2r0W�|��	�^�y]��|CDZ�?L�+�g��a���G�Ih���N�eHx���c�&<���T���^m����Ѡ����*��o	�}�tJEl7{Y��J3�����~�W��#����ȇ��P:O�w�@lz��m�Q6�G�)�W�ת������=��F��U�9�Bx�cѡ���'��h�,��]
r�OD�$�&ܜ�Ǿy�e(����pJ�T�;"�?��'��/o(H�L^�\c���4$mfK;���T���u���hN��*�1D$����hYG_,� ]vAٝ&�IR�;"��Xo&�ڪQ>hxP�邤I;	�T��9޿f�#����~�=�P��NS�ņv���"����CƟf�c�}K�S�0]���k^�+r�	�E���2$��z�T1��)o��I�;AZ`�Zm�8\�{�q���"���K��S?���L�HX�J��-KҀe���^����T����7~7�^��ɐ|��o�%���$�oA.֞A�<��NT��*B��+���������=R�5�aP�F�p5�����N}x���aǥD �EMZ�pb�Tx�Tq���I���u?vak"uGp,o8���˘��5�M7��(c|K��﨧ZtZt�	�xn�Q�Ǻto�1ѿ���#��y7���~���T~���w���/674C-	���a5��l?� f�fM�an���F]�������zd @�:��y#S�~���(y� Gy�A*��HM����D�/[Y��tw<1���
���0G��DJ����dva�<���DB���̎U�H���:���4p5�lxp�a ���-��Pld�����"��g`���v����ui)e[���}ҧ�U��j$+�Co�@Byg��:"`��� �?T�W����?L �kR1]�L�D0�C��ʪ��T���Cd�-��������'��U�݈�O85/r0M4�����h�DU�)��Y�N��l�����muT�.!EpX���OOn����qf���~>}&l��� BN�Oq�\�Z����7Z,��Essk�����QO&6P�DC�f8�������a�B�sNN�Z�&��Cp�T{&��7s�I+�;P���I���Ӿ��f�-2�=���7rܠq�wr�$���dvu̕Ȁ��K�&%P8�Ji�[�|���`����R)��zqf"[�4�ڧ�Ġ�jH>�笭�pȝx�s�S;6�W�C����7Nf�=�M��'�}Ӊ�'��Ο��S-��:&��n���O0��X�c�k=_��<5��	�v�92T��"�RR�ڬ=�?pMa�#��+�(s �f8��Ջ��	޲���i���mju ټ�[��Bޓ��ѷ����]���Q��i���5�A�a�$�?��K`M46��X	m��o�fPy�-�^�d��@̺�uՙ1�MZ���w��nѤD������s<%�bU���?
�F࿠IU�G5���ˊ:��C�����J�4�jN�6$,����Re��7������ڠ�*IUe� �mwB���Z���*ېLj�M��_���8���<�u�9�P��-?͏l��N|�r�/��� �N��wYT��C6|;�O�[�c��Ӝ�"	��d����
y.����q��3�(���6B��Ж�.�%Fpr��{��`�Sm��*�����e�7�l\el��䌭�v:Aby�(=��r!��ϲ$��5�%��e��G�v�9L�ķ���A��#��_m:e�-�N`���k[A>��ﭸ� �W*���a��BG�J��	y"7qQ�,2�}+I�(���?����ø��7߽?�kAy/�q��P��*뤥�
�{���Z�}W�]�����n#�w��,u�47�����Uo1%�J����w6���2���m4�$sQU�;ѕ�6��	���4�� �RD�@l,�<���q�"�%q/�2{*�I�	���zհ��_m�z%�:P�u�I-��F����aZ�s�rm�]~�s6#����(l
�T.�|ʽ���.+��U_氳�ް�>�c�y�����C>z���1�C<�<������Y\g!����^�:�a����L�l��x�;�&`^��T�&b*-<��*ox$�|'��!��F���@K�i@�d,�L��*��LUBr��1g�.�Ó
�o��(RnS�����M���~���������s࿃N��^с��	��"B萎FY�(A�e��C�[�y�U�,�ծ	RV!K辞�ތ�6��@"9�@��Y�Y�s�.|n 
{��CXZ<��-dv�=1#��贕��z��B���Z�� W|��t2<w8�㗙H�;�!��A%ax,,9����f3�z��c���RF���IRǒ�~��8��
C'�@ ��!� 5r=�D~�# =�-%Dىa�r�����O����u�J�r��	�z�����і� �G=
~"�#��蔳����mj�x�p�o����HE�#���|��<�Ѡ`�1y83���Q�(l  �*�h�#�r�V��a�܏���Ͱ���c��R��A#P�z��#�����1{+�~��yb��7���4�K��W)�>���>��Κ�_ە!>7.H��?�nN0�u���a�\l�[����l9�yC�{)�5`eO���+e�E~6�%v��m	�%�i:��CǜBR��$��/�\�1P�W�#�	U��'�[7�<r�1Et��϶/�̽'�E��eвI��!��Wo�J��&�'?��*ט��AO& �{����=9�� D��O%c��X�Bo��J6X�]4���VR���L�1Z�"���H����T:.��Rw�!`�Cp$��C�<��d`$��^���+l(<��ɣ��d"_�a�O�:c/�:��}/��"����\I�$�Ym�$��Rɛ�k{�M�f����{Fǝ�-�W/����\�[�j����pP9>P�ɮ�6�f7��[�,��8�nO����b� ������cZ��=c��W���2~��5�ud�-�5}n��?��@�B3��;m%C����W�z��-|D!�S�$Bm�؆�������kQuU&�[k��Z�?�y���2G���c4���	�BkR_�5�����0�'8�	sh.*v�eLCÊ����@���wIi�s�2��<~�3�_�O�1`r���\~�0�Xq�x\f��6�����f�������PK^?�0��DUhVhN�{����"n�w��j/a&�c��6�;i��U]�ySp�n�u��GL}�������uʴeGf ��e��W�G:M>�m�`��s���y,y ���d���"$LdkI�Y�?,��0r8U�ZR�L4'
�~G<t71����M�N�LǦK����Mw?u򎤺���~g��%i�O�:������N�d� ���O3���9B�f!O󽹜YM��	�E�
衲{0/���ȃť��yKA�qF��M	6o�,�=��7�4縪رF���^�����������'��.ʅμ.�;~�[�g
]��k����t��_�_ЍYx�W�_��E/����袊M�w���fѝ��ΰ�M?��葎gα�\�&y�I%Y�m�����rn��GI'mv����X��0�	��!���x��SzE|�B�O$�I�:[O�%Nr�h��i��˩��]�(�68o �� `f�Ǆ�Q(P��Xp�;�d�)�N_��Т[7�=�ʼ�����\$ZX4"�����X�N�f��45R�!������B�֥=a��!J��tޭ�i�� �v�j����W|�L7���Ɛ2��+�����JX��3���Y�׃6�Rt'�&5�/���0�K��螳�r�~���\��"��eY��E s���Ű��4��m����g�,>�]��*����D��2/���1�N�\�{�'��|�r����m��oM��Lۅ�X@Q�c
V1��UI��^��F�)c�%wdA��1��|>������9jG��`c��p:��&������k���	�w�=�X���V����\qm�����ܹ���]EbƧ�on�4��l_��m-��ā�~�Elq�H�9��zU2����Zc_��܊͟��o�Dm�Q}V|�I�/1�LK���ǀ�i�hk`^ɩ�4kd��dC�[:&�\/H��D���#x�(E�xYmhF�g�礪�*[�>�Fp5|5�I�v���-\�j,��N�e)����1�%Eh.�����5�o����k��%�=����6�Rr���ʎv���"�VU�0i�6kR^����^��B��f��=[[�!�(}G�C*���DO����>]$$߾ۡ��&`j�mrbTwD��^_�C	���� ��3с��T�]�Dh|ɾ�K�k��h�:Z�*O�a�* �����
�ϲk�����Jz�5�OU��=�V���3��3�m7���T��B�\ؤ���9
�w�#�q�~.qu���p>�HJf;�ej0OBA����|�x�-�I�7(]S��V�K�"M	yt�w|g��'D�K��� 
k��~�����}��6��=U�؛_g�L>	�:�M[�����W/a@$���rr M2)�,7齗���1��d߂l�*��p$��e�D쐵���A����� ��~Q�N�T;�ؚ��ؖ���,��vsx��xf`��؝���s�g���X&��Q��$�~�Κ,�팏�YQϊK�*�]���X���T�|)����U�#E���)盘m����s�=/M@n��Z����S�0[W��go�AR���\��-2��'�������\�+����w˜�"�4Y��2NⲼ�U �H�
ǚ!�-�X�3��E��,�w�V�m��,��F��RS|�#l�: n���u�`�?�����s�Ͻq���N��2�L'_02��l����:��y��9M�ۙ&|��q���٣IV����	�[x��n�5>ys�|�V>�s�_�6�|8�K0���t��;�� ?�,��ݢ~C�j��WzϾ����#V\��o	t�S���
G�S�@�9��&�|�<�!��K^u�,������E��H�Ù���<>�hFZE�t]j�0�D���z]�.*�4fи)���>#��)�R��9G�uE���#v{M*�>L�����Z�Sd���Z��K2�bUq����5�L3hVϓd����M�����B4z�.ygt5$��=p��,bq�ܽ�N� ��d�'���	M��?�ܴ J��8��I�Q�g��n,���T�c�I)Pym�����pQ�d:���Y�D��C���S2�����`b��$��i��?�.�R�GIkA�Q�U�^�n�?�LU���}ǹ���/�U���M5/�1Uڥ�ʑ,Ψ��f5{�^Ll�`���0��+L�/g�� 0,��>�\��p�<v�pe� ���*����_��A�QiH��O��iK�����X�߄��Z�F��a/N�/���.�ZD��$�mJ ���4������%�z��d}sʶ��'������'�щ�!5�t.��7@��&�����KI�����8Ǔ���+��O��F���;x��4HM���y��4��#B�lt�����ߌga'G��[m�%����]A���|��9i����ǔ@fB��vF��}��ؾ�Z�a��#G�`�Г�2�z�{��u�(/R��(���)
i0/f��@�*�d�۠����$����`��m�?%�v0��/ގ>���d�`�t�ur�;��4nг��q�d��3��3����d�|q�����P#O.�3킥v]��@V��*jy|�s/��X��_:6`X�~�m�Z.�Hh;��6iYzL��͹��n'�K�����}A�f�o��g����m���J�ӞT�`�	j!�f��D�Ȼ��+HS���4�TZ�pz"w>jZ�L%��J<��=.I�;o�hv�a��Ov~���e[��X�xUL�@�V�F�<�s�|����Ah)��ok+�N$�5R����~�x�R��:F
��x	�m� hq} ̠f`�3{)B[�l��zOo1�-á�&�r+C������g��p�Difg���+�Pƃn��s�f��8�ӊ�R�@��ִѶ��j���~�����F���PS��6�^���f?4e�a����}�2���!�x�?��_HTV�TO�B嫡�}8��x�Yf����P_���T���N�4.�:!�DYȅ�������6���u�ӱ�jH� b �v�`�@����.�G���
�����5�iN`$�֋z�	����[M͋����{�=���1���$*�3|ֽ?o��?���l��e9W�2���?�٠�G��;���grZ��k�^ACP1h�э��uV��h�/��2��{�����v4?	d�7w㿧�#�E�ⴙUd�E�N�i��=z�9`�|5˂�
�76�Q}���4lc���"����f�H�|5W�����ߗc���ӔG.��HC�,���L��+a��7�H\O����if�����c0Qd�\��g�T:G�M�	/U�\�7�wE�qG��������/ψOUn����_gLB���4q$�7�`?��.���I�"�.��e�֥����Ȁ_d�ޤ�gҼ`��1�%w�?_�J�Lo����5Cf�L�K�+�&Rh�/6M����u�z]��E Z���a\
�<��+ٛ�6�Q����3�w{� �{LMEW$ݛ1�ͦ��]3q��l
�8i��݇⻏(`I��؞�w�Z�r"����cV�ƥ���`J��B�̤a�Y���b�f�@�m\�n#�	5�_�q@q ���}�v�lAF�zh�R+��{C�*z��["&�ِ�*.�X1��c��3�����^K����yğ�w�����~�2�0��$V��٤�ri4�RMi�rBy��S��3#~oο�>zՂ1���]��:cu�\������eC^:��9Q��O�P:y�6�B�ͺ����|x�$HK�=������:�
�_��P���Y���~V��-#l�r���E`u������j�i3��լ��włH���F	y��U2���K���?J�s�����C�8� :1��7)A�ʽx�G��[D{����lz�HbycV��ʊv3n�]ϛ.X*s�f���If��lV�����b�Ig���8�S��\���������/23f��na'�|�+;����ѓ���꒨�Kw�w�wZ�p΅�9с�՝�u���6{*��Y�̉ �uq*�K��Q0������m?�'̿��*��H�![�t�s����`��/g���.�[Ad�-0��w�'���"v]㦻~{0�4.T��ǆx+�=M��f%�g�o䠈T�
��A����� 0y�\4�&Q*���C�b��1����&E���*�g` _5��Q�Rp���HS^��V���on;���^��8M��f�s��'c��[���ۘ�QU�x����۳P������l�{v@!�Տ+�Y�?e���y�)�ⰵt�f8S\���dw�������-J S��`W;E�D�Xc�.��⩄r��sg���
���!�G-j���ĩ�\��J4�zӧQq���v<MȲ�x���9SV ���5�Bu�g'��\�YG�'K�z�)�hӔa-�6�9�Mq�GCн�},��������	�\wi-�4�u�cT ��0��~Y�r�I�!s����g�L���E4` �I�G���ĸ��㘜j�L��9�sܹW���<��W�ۤ����.���K��8�'���i�N�u�D�����-A-��8)�<���.�+���vX��Qڙ� �m�ӄ�C�-���=�������Y9|?��$�5��5�w۠m�˨Pz����������V����β�o���#Q{���Z٤�o�y�}�9p�ȇp`^Ʋ�;��K��S~�����9�W�}x�3�?.RR�
^'�\�����o��chB�2������kZ�sD�ၵ�t7���P�����"w� �]y��B}�A�VH��6CD�ȱ�OJ�'जa�NK���j�[��(:"i
��Ն����n����4"�M��7a�+Ǡ��0޽�
R9���z߰K!�2Frȗ�躗��hM ��j�o�[)���ݡ���wq��ʷ�Lv�E����&@SyI���."Ǩ�8�hC�&�.��o���\�ut��K���� U�p���gA��L�z����h[���9/���H��W<�Ĺ3�\���(�,�쁑�p.2�c��H�v�>��mN�]��>��%��&��`t�;CR��ړA��ڸH��~��Y�G(p���ѵ��9��( ik+p��y8|j��s�^�c�[����*xY/�颥M�HL<�s�%���"�7ӫ���gq®ZN�q٭2��$�_�.��i�p�y�Wh��$�y\�eǘ5Y3S�-�ivk�}��;-Җ��~[j�˟ʕK�)59�ז�R����Wou��_��i�2zA��{x��H��¥� ��ޯ��+������H=�fp&��2�6L��(7sJ�^�����ڡ5p�9� �I�YP�
O���V�eE&99��`����
%ا������ή�Uc�����,ɲ̽����ۚ�n}�q�r���J��c%+��MF�pr�84����\�d�O�-vmК�a�x�0H\�� �կ8��v<�*�A�̍�����.�(����	')@e�o;���7n_�˶FW�a����v��Ϝ�Ǻ�_
���7�_$𤾝=��� #bړ���Zk?�]";���[z�.T��<䉃3BY��k�SHySPc�����)��V�7����b���B%�g��^(w�4��;���v�T��ʚi﬌c��� ���:��[<�yh?c���!x!��c��fJ�9A�{��U�2��P��R'G�~"q�9�HX��n&T~o���ڎ���4JgO�����ܕ/�\$<�Iӕ��d�p���Vt�4G��)ż��8$9Seƅ/<"_����3J���H�����N�4���@�,������1����Uk|45�;P�76R�è[B���RR�����P��'s��W	�j���ELv̘��j���iKP����T�=�=��<���,+'*eN�	�>�c��G����fI�W�M4x��]O+�K00�)+	�ӂV�s��'���GD���1!?o��t�r[,O�6g���s�<���]�������5���"ui�IQ�`����]��&�zF��N��V��t�ZTb(;cB���M�l�/���e |�ۇ�];�-3�	
9U.Ny�n�֫D�%~q�x�/�)���^���|���`3��,��	d��<ɨ>! s�T�1���ipͰѣN����ŗ#q��R=<�n���ޅ�:�vb��k+�>��S��ͫ]Qg�m����h�)�0�ǹ���JW���j� ~��[�{+3Yۄ�z�*O	������M�� ����AB�h��6�R�\yQ�p�������C`1|4y�DP ��iK�z�m�cųg��A�4��;]����LK������Ȝ>�g���6&}v�'Ò�vle��礚7{_��3]����%��ķ������\LS����NRE\���񨊁�F�O���j�d�P�ޱc����w3���ຩΆ�����{8��Y� ����]��cBO�{
�0���kw/[��z���N�G�9�Q���[h�����j�4J� ������"����|ϐ����οK��r���噓�xA� i4i��5�m:F��l�����P�Y�+�K�y>6 W��+`B�O�����Y����%������Ͳ�P�>d�����g:%r���xm�]@��L�����f��u	�}�no�*��K�Mƌ�%�yq����&���jn�R? ی���K�S��&�����-�t�����&�%�K)��6\���`��J�/{�N�P��������Vʡ�|�����������/�&���K�.y��+ һ��g]E�`�j����e/Kg}���Ld��y�E�����1���v�ל�B:a�1X���w�:��(};�,d5�K���,<��2ֻg�7��<�M* _7oW�z��vJH���`<�j4>���ז0钁���(k�y��3�XA�į;�a��<`���`�υӭv���Ӫ_�좭%�ڇC e���2��T,�$ � 0�;���G�I�����xSp����/UD�;w΋�&VjI�����+���Fs���~s6�m>P�����`�;�֑Abu�bY;mS���a#\;v�Q�r!��}��KG�����8�$��o��s���s��Ö�1�Ҩ�?e����꣤�q8$Y^i������"�l���F0@#ȑBLb�5B.�����2�M�m��r�����?JA27��}�-hLS�ۂ�)(�<c\�6N}��L����LlD̉F`{�B��T�NZ�l4W��yr:9D��v�ȩR���dG㯥e�5ӝc�{�ȕ|*��7x/��Y�:`B��ˣ-S��2M�/I��[�����#��|�׃q9�
��w���ȗ{�;���'L�*b0�;r&&�<{�2YP��
��G�k��B��e�����c'����j`;�j�eV(�1O��m�����;���K�G&���8��t;�Ϡ�N��)��6�h5txl����JŬ�(���9Q�9��?�
��)��nuCe�P+a���6�IEhj��ihr	ä*���Ε<�;rS�e���A!��#g��*DV}���~˒fk��q��,���1:iSiO?�U$�+�F�y���g�h�p�)t���(��L�d�I�	"�K���YGl���9R���7XU��]�F�a�n�����Yy�_�e��)omalS�:��W�I ������	�`0=�Kj��鑱��nmC�Aj���b�d�EAU���v�B9H�Rplo<E��&3~Kv�*P~��u�׌�8��K/ �
��]��஫�s��AԡRz}Kз�U�, �Ӕ>YF^�l2K��b�)����
^��E2�ڜ�M��E�R�N�iˀ���
��,��ݡ=�ĺ���?��])<BL�^����l�ey�&6�$�߬rҳ��z�K+-����s�!���9��l�'�]���@γوV�6��p�M��V�#�#\�d��rEK���
���P�\(�R�zv�~�2�~�KZ�+w��u�l:�D\}8_�����#P9����DZ��n��o�*���"��be�ꖡ	���v/w����)w����J�rGTv?���w־���U�g��*�%�q�G��d��r�����0��s��4l Й^6���H�E�������v��k!$r 0*����	[���{p��QP�?��S{�[�^樺+2r�ldۮ/Y�L}[Zs3%�t��_%\�_�= �	ol��.��,�y��۱w��q>;�zP/�g���o�J����d��-�/���`*����|(o�V��L(=7�!x��	#,VI�_g��d0���q	���}�'ޥ�+��!V�}�>�4?Z�@��C[���U=�q�=��:���������˵�G/�뮲�79����Wx���Ln��ɚK�����:P��2+ZwG ��o��W�{+6��r�+����D"�<���+3�
w�qy
�_�V�	�oU�3����7�Yn�g�z)�uљF��������R��Y�snu�Wkx�*PypR(%������>F����#r$�S1���za���4Wn�,;�ƭ(.�M����H��EI2l���P>
��9�x�}��#���O�Z�����x�G��&R�6���2%,T���A��^�Qұ�m�A��z�S���;,�*l0��~m
L2pw��`�a�A���o3u�e�X>���%_UL��n�L��6�"��c��)����6PԴjb1GlBi9�A�v���j���͑E�yO��G�׹�MP!?�eH2��	��h��`B�A{��^�jo������%p�1�Ғr��R�> 2vbe	~���O��c,v3#�5V�17�_x�뽱�Z��v�]�N���K͜#ᅧ�)=��<��Φ�>���.c���ܪ���ɵ��3??^�k��b��o/&_D��R|g=M\&`!��q����W�n�t��';�*a�}H�=�X��Wrs���R��i
�(����#��0����pc�Ў���%�[��N�c*�� *t鿪_�q��o�s�:H�#�̨�җ�4��SR������]Qb�I��*Cq��|,�n�c����C���@�� t�������y[t,��d�����YILC�ު��1č�]���,�]�0�6�����Z~k�%-M�~d������/�[~��)&0k��W�Y�h�`UεDb 	��#|kX�h�+&%0�H�����N��V�"�Ff���Oi���W���iy�<Fr�	M.�^ͨ���`�s/P��R���a��<W���M���2����{+�@�q�@l,N˪x�*�jP���D��.JH��iFE�"�ȼ�)y�3���G���ӡ{���=��db�ܑWs�I`�g��ˈ؉���y�]���O�R��q�-�����ەP�p���L܇����@=	�}�y�cW�b�o��_�M)�e��aK�~���7}��p�1h�y�7Zȫ����ٿ��+_b�n~"w<ϕI52f��d�< w|(w��|y� /op;Ej��&�)�+�����5cA�
�'@�h������Y��Vfa8��|U��Vt$���׭�J��D"��P���h���rxb��HA .���`R������XE��Cp��(��*5X�GZ;�ǎ�8-A~;���V�}�����2����lI���!���A�=��̝4��`��7�m���[7�?��NNy�@Z���s�%X%S;��s��U�`��+QUL�i�;��{�k�!�U\��AR �v%����7���IC���!�#���a2��P��U�lBH�Z��[����7Y"Wޯ���kͿ�4Mo�t�:�h%\���R��K;%O�n��?[�C�Z�RC�@�t�n�8,;� 2��k��m�����tM�Y�1������$���_��/e!<���~�v�iEE�>R�N��;(�J�Ж,�����j�e�~Uֻw�<�������yB]�7��nh�ĊZ)�u�r�T;Ё�*'y��M�������u$���s���CZ&���4t�n��U������x�g�H:���a��,�{��P̧]�wd+�(�=�f��� ��I�Ԋ�*N����u� a����u����X ;�.��'������d=��l`t��p�kW�C���Zc�E�5��)�xS?_y�t	,M�@�靺"ح�~�홦�ѕ����,���W$��s1�+���dF��8��/Uk�K]�1�&T/Uk��]d�aijM^�ԝ<Х[�7b���=<z��:�u��RƧ^$���R[;I�t��������g�XV#]i��-�U1�B�s﯍\�syr+��u;���S���4�Է[��g�F�OY~
���Kn���P��s�s�7U{p[O ���hM8x����L:��>u��|˕i�`��UDZ�����tN��K7��e=� �V���zAC�3^�1\����=a(�h�)����	S��u}��"�˓1�� �a�����w�0�n�oFa|`� O�h()
�&���:L�hw����4�Tm �� P@*��Q?-2|v����o�h)��&N��Y`�ÓԜ��A��V������������7L�M �>4��S��K'�H���]L��|�օ���H傑�1܋np+�!�LQ�6�`\���JE1ٓǥH��NI6���DE(�
�Qŕ�~���R�긨䑱蝔�ȢcO�h�[ɞS��2hx�w�`jj����K�׈��=�x�~�q���x�24�v����MD��� i�be	�i� i����?�&���x'Z���ؒ�csn�����Da�4y����h�|N�����6�����Iy&4Q3��xr�wI��y��=��0 `w��ìk����41��h�O�>��tD��)�B��2i�c����R/u�q�Dw��tF�S�l�_�
Y�^�p��wp%CWj�C�2I�|K:�v��'{}�=:fԙoQV�7u9/��ڝ��&���i�-}tY`�y+��4�7�8g�kK�q�� 6M��S�#���Mg���Խ~���!�}������K��S1s[��`;�De��GC��;��V���y�������=OZ1q-��5���T>�ybʬ>�1Wv&Iv^z����a	��g|�8��_��L'M�w����Ȥ�v>�?C{���S6���X��ߴ��OΟ镒���y:���P� Y�>�C�6[ IȖV?&����O@I����q�8�n��,E��2�2%�Qm%�/r�г~"��������8lJhX�p.�x�dA�֥Œ��̣�o�ǪA<�,�|�x�׋�u��#G�X�A�cM���j�l�> S�O/g��[��P$ǔ���f������?~�u�y�i� �Gc�&�^=8b͉	w�ƙp����!���Ԇ2�-���?�8��L�q?��H:����ʼ�{0U\�'4��I��;9���*��w�v�a���Yҹ�	b���p>HOū�v����?Yͺ� �%��V��M����(���4q��}T���|������\?�H=����ѯ#\A���롩�q�{� ��C�D�=�Iw��U�����m)����G�C_il�ڋࠉ9@�_����.1���I���R�-/���}���>#��:��2}A�M��7ek$'��vqHH?��$�|`���/Kc��F�F����(Ja�f�>����~v�v����v/#�q-[���7�����M���b9�D}��Ԭkh�5�g� ��ހ�{�2��u?SE���
ˏ^Y�~��#~}�)�W���xiѵI�%�;�Sp�J<�F	9^�_�%����6�P��[»m��} mg��b&J���A^7Q,_��r~���BT��	�����>{����n��ێ�ȡ8��gB8T�R��!�l=�-��w	F~V*���\���{ٶ ��Ȥ߷�^߁{؄;k�[-:����>�/�Ic�d�1��yQӓs�� zՀ+P���v�3&r�a���\��aD�!AFBy����,��NH���(h�)1���Y#FNh�zb��ǧ�Ώ�M(����(i�$��y��'W���9�1E�⿾ۦ�ŋq�<�1���@��@��OiMm=m��v�?��G4���^A�}��X.q��dD�I�8���X�HE/�)ܡj޿ʸ�0�sJ99H9鵊+F�ז�G>�:\2*�Zj1>ǔA�����ɭ^M-3&��1 �ޠoh"�x �����G���`!.=����q�|v�����0��T��Cz`j,>)r��^����tm۲K��]�34�����g,H�� 0�\U���g�矫^R�P/9^��4܋JᚼT��[S0X��_����6>��);��S��y�G��gm��|�8it��ę��_����S�<���A��cd$iq��[�l�;�f�p�Z[P�ju#s�����=֎
�t�G ۆ@��{=O�C cG��R�8(����WE��Y.��i1�c��*����[�{�L��(�Ag��� ��	I:9�v�:��x�Q���ۄ(��U/M^�(:����t*��q��Ϯ�a0Z=�c���t�1W10a��P�I6�2 c<�+<�9
[B+�y6��^���w���M=�M�f���oH��S��ԍB$��׾�"�y�TH��A$I��3c��H�Z��5cs�٣���L	�	82� SU��ML1�E��>�x�ռN̼�����$���6����~vQh�V��B&�.O�e�����-E^�ͬ�qhX����>��:ؼ�@�tw|U�ٖ
H������˻z�� �c�°�WdcIGo��(���)}+u���A������C��j��gt��8����L�Zh�x��2|��4W��O|8���d���p��Kx���h�a��^����]��'��X�w�n��r$�A|��P�ՌS8�8I �dJ�"@����7�GY��q� mU."C��}t����n�.��\VV���K���Q�(kKi���y�q�u���g�Ӄ���vL�۱�x�����+*�O�H6�c������ZY��;�bV���p_�-,���'��E��Vj���✽�x��\�'G�\չ]�L��[�O���h�FxY�Ho��9�o0�`K��~�S/�`;�с��9I j����]M�}{�ɷ'Ă�H0`���	Q��ϔ5��{�2��]�y�y��w��E:�7���S9��Y  �N�lA��4��zp\I��il|~��]���2������te�,y�9�^x�'!�O���Q:D�9�z��p���
�� ��/(ȟ�!zB\)���j�Ob��O��ْm��ޡ�����"?����q�u�C���n��x{Y�r��l<��@�]��4rX��_��Pփ#.���aOK +(8��jY���2шˡK���_�h�����N:#pR[k�bnXӐ����a�W�yM��U| ��Ǧ {��9�&1@�7��X�i�7��oY��/{��Y�ĳ���f�sdHN"��.��B*����e�}'���+=a̓�~P�#��
=���I×_�hJ�3�p��a��
 DR�f�`3)b���{u���$�!����%�e�| ��?���G���Ų��y�8	�[����k�O?��&�������u��ئ% ���}��#���t��Pu����[�h�}�$�.d��B'�Fz��d���?����M���zC(�tf>-��O�Kw��S�H73q|���;?R.��[4�T�t���+ ˖�y]�j`�Ž�������Ug	B��z�x�����P��t'���P�S��5�O�/�d��H�V��ZW
0����_��|��@0�iXy��a����L�<��*<��=0B��Eʜ/��q~�;��*F��J�[[��|��S���5�񒋙�^�p��Z��եX�_�Ȃ��WЍ�V@AG���6��3�%M*�f¼-.���T��3H����N�'t���4�5��\���e!t]I��hat>�SR���TӭO�w-f:d��R�a�D�؂߸����o�)Da�(����vf������3X���^e�jq������t�H�ش�ɳ+�ĭ]�Tbf�E��6s.q0v)"���=��~'4<��CG�z�/�5)��c����ry���V3��=� �r�����,py�Z�s���e��.�?FFbs˪�����TZ��W����X�gc.[n1�Q�g`�H�|�����]Z��W�� ����8 ���CK\�A%�Z�ar�4�[e�y�!��-{+3�?�=��"�#�D����P`�6�2Sb���T��V8����3��v�D��a'�+�U#ƿa����Gr�D����kC�y7��m{�f�)�p�Q
·oR�Q� {��)2�k�H��o�(y"U�8i�7��苐E����
�YGp���4�eԈ�p�t�صD�9A�A�?;�LM����З�{l��r�:-2j}##Y]��7�,E�?�r��Z��M��q�)sΏ?b9�X��U ��g���`C�$�l�J�W��.��-����[���L4���QƵ�:/�%k�L>1��6oBB'G�F�g�dp4]���}G����96�fi�-
ǡ��/~��4?�ٞ�Q~��F�-�n�`�IM�a���a^.�C�O\�D��eHmԳU�0������y���7~6J�G��a80֟�f��p\s�rOb�:�f�.�DɅ������&�#r]�.fFS���h�:��Lf%X��5��Q�r�����e7��?��PW40�>��Q�1�uJ �j����b�A�\ֳ�d���>T����0ʿ����G+c4�9�� <]���0g�6����U�Zݖt��N�w�ir�;�>t��/ٜ�0�\>���LƒsIA�d���E
Db����W`'��3w�����dB�ˈZT�ls��.o�#�`^Ӈ<W�^�{w{��ILT;n\���P��Ά�G�O��eشѧ��{C���A�n[Y+d&��m��v�Y�%�
����t&L�+L�L3H���m����0˨(�Qn�66�ْ�X�q3���, }si)c)J�1�w�ub4��W�#	�3KDS���,�buh�Y��o���t�\Arί�"���g�W���ep(4�&U��6K}E�@�a�D,�}��l^������Si^�AHmVQЍU=�pʡ���W�-Kg8�ly, ��w��f�ۓ2j��)ే�}he�0|�=P��Ǚɯ_E	���ΣZ��ޑ9��M=�f����?�e&����\��q� ĚʂYǇ7�B��(�'S�ԉ���Ybd{����/EsyN�!��}��dW_2�����>$����y϶�]/ XT��AϺLZv��hWa��D��B$�*���|�( ���ˠ����6��g4C�9��U^�"����V�E|��j����c�a2;=U=s���� �R^�֔cM��iP��v"��
b�;�V��>�&�b��	�ǡ����m��K��2o�7�ZLUT�����+�<���a`���T�g�r�Y����7<K�r��i4�9���ͩR���'�
�Q x��7����:���y�C�\p���wӅ_Q����o��O��(i���N�"w���>au��[M�Y� I�p�ӆ�C�72��̙�V�m�j����.I1(��T$f��`�o_�S:B�� ����@;���/M-Ŝ*jP_��3��t�J�kشg�!�zm�h�*S�z�Et�Q��r��n�C"�Z�;����.N�6#b�";*���T:�<b?�Z�X�?��[GO��<��+��o1\kVuc=v��m��-^B�4+��$�)���L�:Oڥ�/u��L��)��!V��?�u}J�a��E�q1C����F�ya�E��m틺Q���\H���g�7��Qx�ol+�CRb>S��u �V�w>��I�?1Zr/�X�3�P��z��Y[Z��ƹ�V�c<�ll6�\}����28ѐ��x�'���_����|�*&���:D\�cJ�i�������"Y����p�~����&�d���P#�0��H�Ď���	Sf�d�t*�4�p����'�0(�I����z{u5�<�jA����1�O��ґ��)�X�Y(qF	TT#(���ZqdL�����X!�L%�RŸ��7�Ҷa�e���hN�1�};bU_?��Y�?e���b,i\nP�'���@�A����m����ҵ���*sD��w��|x\�w��՚
l�̄�÷���e��L�;�ɹ�7�qbr3X=��Wn��FH��pܵ����V`��]�I6�1� t=Kn�m��~�J�3{LF����
Bpp�B��=0;��q�,�)��g	�/&���	w(��
3b�d �*A.�"�aڨb�,���p��-��>�9U��w�K�,�P�*�Sbd�*�b�����P̰sJ�[/(�qH��S"/�7����=�Pp�#�!�ո���J&�n��f�(j<��wzo�4b�Z�6ຩ?v�f�%��^ڝr̠���Wj �w��ȋ_SRo(�c��B���Xi耬5�(kS�Na&I/�n_˄ԓ�2ZC��׳��L�o��vZ�V�a@���-���+�x�7F��F��zP��,�����o4��İ̣,`�Ǭ�}�)}��YZ�b��"\�ۈ�Բ-�m��7N:��F`۾�^��En�������C�o�y4�\��uY�R��&,�{�pN���΁��8�(I�j$so�ܝ�f9��`���Čƛ$Ԋ��n��3��z��W GQ�)�(���&9��Č������)Ȍ�5>Ca�~�ЉA�C��AcS�[	�p��Qm%�5�0��)��W���7���ݹ����Y͡k���li��b�o�^�����]}���	w�;�isl��{�Xz�,���%� ���������6�M,<N��`��:�|~�� ��������	 ����ЯV�e�����[b�^+,��?�L,��hk��l� 2%/g�_��3� AA��]�bI��NTbY���{�m24�6��*D������O�7�·�_���@�CʄB!���7(�X����[š���<�	(H�������n��4����gz����Q��)���E�M�y4#���9��j�-�pw���V�#��$E�8�8��7l_�mM�u]���@x �%޺̯S�g�:�.:��Ա����~�zd��T�Vwq����a��i��:�^�%��<�rS��Es���E�ڢ����sl(ǋJ�����̄��kE��9"���6b$4���Au[�hɔ�@�����?�L�i��Ɣ*�����*٠!ơ#����<���^�y(��⏇@��m�<3po��E��������w���-\����V���������E����	��ϐ��P�_1��J�f�7���;nդد'ɭ7
Z���S�� ������r�JH0?Օ��%����Q��ŶD��~j7�&;�v��3��R\`b���0ݻ
n�|��m�yFt��@&���qx�҅u��~Oe���>Ll�4�X0��B�Wo��
�%�#__���8%��c�t_�lb�TZ��*�͒�G� d�3��{kM�@������A���+��۸v.��p}�"�[�r�W�R��h���"������ck��C��sU�m��dax��|f&��"֟*^Gd�M�Am�&l�E��Q_��(�c�ͬv��c�ۛ`�RI��OY*��zZ.(xFZSM���Wm��\-ɿLF���x�k��8M�;���O����B��XJ�q��VdWp���$��v�}�ʉa�a����"�U�b���H�K�Y�/��my�"�TF� ��H�K��ˉ�j_=;aM83~��zx��]S,��O���J�p�l^'���:�t����;��3����sͱpɊ�5\�JjLHq�$�	��pa��(M��2t�L�$a���k��Jp�j���M�ooD���BX�S�a�}+A/{Dw�C�E\�!��۶������.i�5���ȱ.�D�$"�$||��DJ,V�aQ���L���Zp|�A~#�g�VMt?X+�jO���1��{!<��h��]c�H�=/���>	'�*���l���ɝ������v�ݗ�s��yޕM���N�`�Щ�I�� Vۧ�{�lD��o��͗,PFp��Ę��kJ#�}LSSه��T~�m�\�ts���++�4n���^;i�tW�,%���w�?�gŅ�rg��nmO�K|����Z �U6��֥{����I9�!z�RG:��B�E��������_��A��FW��_���e�('#'���K"�sҫ��VЌ+3s<�E���Hkq�F�x27rn���5V1�0�_�v��H��?��ϕ1���Rm�qǭ0LI�4�^��KS�^X��p�W�u9�P`���`�N�������3�߾WБF*���
�>t^�>3��xj�d	m�{=X�u����ߓ-��/��? �F�<���v%A��P���w肐�?uU��qB��/�LǜG�����d��G�m�Pc���լ4�գ�
�X�E�j�� ��/�e;&˦�����j1#�G�s�Ӻ��*�0�?�|x,P�p����j-���m�b>��9��D�u�����Ԩxg`��a����\q(�Z�z��B`,S!�TC�Id�r��)jN�x%%�y�.ҥey�T�����dkjf":�W�	Ft9�ac�y�V�ܣ�v�rk��jo�����o�L�S�����/�K�4[����%�>��Y�p���
��i��A�����p�뛳Ӫ���)B|wM�q�6D���v6�ʛ}~��r����.=��F��{a�)�|'�/�4�Pxѭ_��l�N�aX��1L���o�C���>��*KfI7_���R4hU�9lnv�:�y��!��wM*i�	qo6��C����g�O�x�i�9��f�Mp�͟蔹�"���'�Om:h~"Z}���w^"��sN�)�?���!��� ��2���=ϊ$"M����?��*���ݫ[��~�=uq�t��7�����N�E;Tu��4��T]]�Ɩr1��(#[
歴�"\��WF�L���b�\���&?�{eA$nkr��Wi�%iB�#��5ŁW;V�V����X��:/s����42���Bޙ%�T-v�L�X���ǔ9h���Z�9�ƃ���Y~CY�QA��vP�?�s� ���8>{����y�DI����<�m�"9�W�G��t�ӭ�Eqp����F�@�^](y�L�Y�`�#<K*���q�?
N�(,�Yb����V�3?�;��'V�h<��@��MT
�s��>��Cu����b	�l�Zf)7�u)\��ZǺ��N�	̔'�I�̍�>tv�s+C	���6	�#����Ko�&Q�yt�-���Hr�g��!~�d%��!?������m��%�.���'/�n-,0߆՛���cE��XPDܵ��H]�5�Θ�C6�[
���)/mlU�ep�m�L��n;$�9�x��'c;�&ț�t��6B\d�#FZ,��^(�̽Z�z��O(��=0Y_�rx�s������v����"�EL|N�D����s����8h��yf�l�?K_2L
���YP����-��gӕg���po*��Ѷq�e$.�8�1e�S^�>iE��f*B-B �!���Lcܞ|�ž�=K�v:�e)�1�N�-�9��j�i����z��h
�:}1�X?Ր-���
��<���v+N$�O{;�]��Hsm�4��ӭ)%�Xs�@������8Ռ�܊̗.�z>�Q7y��[���eH�2��UMF�������D�nZ�n'���c�
uF=Ի  �tJ���.,��o��.����G���0{�����:)�@.���"�r�>*�y��(�?v���U��!��tn:��^�܉oO&P�D���x��N\�������7���³��ކf��u�W5�P�=m[Hh�Q��-���
���bi�p���c�[����:�}�$�� ]2ej�J�5��e�k<�Áe�ֱOQ���[ߐ�jJ4KǱ�i�<>��ꖜ1͉�8u����Q%ȗu|>R	��`���1�^J��S��غ�Q1���M6N�#�!�-�J4l���%��p���2�`fW-&�О���n��.��AQ=�~�u�Yg�ع �5�S��ӬqS�5 �f�x��p���
�YzT�۷�������燁Ǟߛ+�b4�qq14��@S�2~�rb�GP,�~c�����1"��rPY-��V��LsԹ��I�<�83v�F����-�A�1�܏�m���5(�ԑ��3)�L��L�xK8��#����Hx�~���sKl���0�o5�v2�����wL4M�(�LzN!4�N��C��DEwv��9"��s�ϩ��\�y��\�
T�Q�� ��oc��v�>c&$~y�D��Ol�3X5tm�}��^<�d�
��JJ��Z&���.��or�����dLp�ڭՑ�f�@h��C�ȱ��3��*�Y�������Ic4��r9	S��6b���p���A�)��0��2��mn�Z�ξ���:��*���9�\UT~�Q"z17ڣߓ��
�c�<��v�݌�I�3���ԣ�,"�a��R���5� 79o���ԲH�"�r��д��7�;�Gk73��<q��M�Ze���;=҄�Bq*��,X�k�	=r��Q_4	�>�ĭ��l �bSP�л�t��r���0N 1�駤��v��{}ϔ� i��ܜ�����Q3;7-?*�ai�r<�[t����jU�9R���(Y0a�;�s�(&2z#��)�g� @���ң�zW�?JQ3ՅC#L�;�Ώi��4^Sh9��>�ؾ��~؆g?�C����"-1�W��,�$H�xǥ�_x#j5�J��&X�oVz"��p ��A��?y\����w!�+�DM#��Y4��6���pT_d�!]m�U4��bF�Y$)��e�����"�W�ݐ�
��Ά|��7i�'��P�}ϳp��S)�z)��5�է�k��jwe�T�v?�����m�W:`�-;c�oI�?�W_�.��.k�W4��rb����d�Ӹ�B߂��s��:��FN��ތ��?M������nC-�e�n�=찔�M=���鬅P��G�x����Z�h�$C��	��a�;�e4��Ն
������	�V��>�Y�����q�d�_��$��]���*R&"�Z��>p�u�w���d�����<���8d6�͕�4\6DE^�{���{N�{w�i@D&�%���Q���1U�s)� g$��v�j�n>�D�7SO�P�n�n��}����M����'���\LYkJ��]�Ӵ���ՙ���F����Hi�h����nLg	*6�2�/Ff���f_��0>�~�Rg�l�w9�����V�k���E��ۥ�1���I.�l;��^\��T	A'��S�e�b�E�`������x�o岘���Q���3h����[~�я���)/���iW_2�5p�=��?}�)����O�9�	8HzK�A�P�i�����㴔�x��,�R�W���#6��h���_�)_py�������#�3=J/
�y��K*Ԩ��l���/�����--�1m�9�Z��^;9��ȓ�Y�-�Z%`�P��_Nw�V[>a8��zVT��2"�:�F�JF ���#-�hs/��7,D�.����wUϥ�u w/��&��Z�ZW[���h\��q���?�ʽ��  �9?����#�/`���72�y̹��g�����E䒤�K}���- �^=��q���(�sf`۶��Y���D��� i�o×"��,�T ��<�}G��3r�v���~�<(�~���o�b��H����F!��	����x2|}���ʊn��1��R��F�Kz�d�ޜ����sʂ���wĝn������!��=��L[����"�-����v��rV�L�����G�iRи�s��d��)N�F�nkI���a�P��$�[��n
�y����.6V)�;�����Z%������)!��+PX<��*���2\.��GBW�o�uOϦ_�@wnt�j6@��5ZA�C�}&]Cn�ķ|��k�P���d����}���eYy2ఖL;Ɛ���8#�8���ɿU�X�TF����?����
��c�:�͝��s).�O7�^��S�(�S��ߣ}��'��=�A�}q��1���"k(-XBȩ�v��X�M�3uB�b�
B��5�d/�������9�T1"�~ڎw8,���e&WoEY�u��w���+$+bI����Bu�c�mY^PD�*�gn�>���Gb�\�e�S�1ǚ4�6�/��M��������'/H��f�龖R9��`�4Z����x=�0�x��V'��у�d�v���i���pC?��6��Ol���G<�~9z�s��utf<eL����
��[G?.��M��ոi��0��՘lЬY����T��푯�~�)�*t�D��,�Q��Z�9ǥʴCqGt�	1�̹�o?&�\Zw��&����B�'"'�az�e'95���B۞�~J��΍�&����}���'��=��1��{��َ4��E��iS6�j]	IH/�f�Պ*��a�;wU����\i��Z�}7e��!�F=����M�5�YF׳S:z5y.���:�n�ŝ{)�DW[,ix�K���]��/�1K�M�W����h�nQ�65�V�%�30}�0	)*ؠ����l��%������Ж鈩�X�4��")�eC�Oj�1ɔ%��G�J4�*�����u���G�S��p���N��-�Zl��\.J�3,��_��89�eYZK�u0@�_~�7�<���0K��_�b�<��l}p�i��m��G�_��d�3��@�#΂�=��e�zwm�zw �����X��(c��>5��Oc��i��L;%?L�M�!���u�Vz�t8`��.�*Ω2�Z���f
e/T�'�i8�*�[�Qy�R������v��Fz˽B|��f&�!W�xN*�:�Wg�$��H醠�Z)C�^Qrc����=���R��2�b�g��
�f�R776���}>�4©nA��( 9��E�ِ���&<M�x�⠠n�1�#��%�q�	SD�G~%=:qzc�����B���k`!�H�Wֱ����?�۬��Zi4�������\ň�Ό��'	4,|o*�p�
�m�;���iz�������~�ar���sDt���cz�=�c� �H���X[}�3�!��@ꋀ���	K���[=��q���B���9%T��R�+I2�z�,>������2f�p���/]�^�U&��w#�5r�qEv���QkQ���;� �T&��Ͻ�P2�B�%��e"�a�b]m����U�)��*���I	��x��������\hᡝ�������3$�us�H�7�\�b�/�ԏ��Z/�
�0c�*�S�3�!��-�|�2�f�k��;dB�k�� �QBD�r�͈4w���ާp9-`D�_�!�V.��Ƥ�"�ST��P�zLK�^Sf�j�$�qy�0n,\�=�����";��MSc�G-J� >ށۗJ�7����{�[)B+U]��������PZ�r �8a;�'���?+�	`.�{��#�#">�s�O�Ҟ�ƈ;�F� ���֣TnN+��@�atWDe��j��D���9�J�+Ueh �����/���r��Ӱ&1��'����QtR^����Z����B<L8�b�,=�N`�!+7��\����f�`U��![�4<�E���l�nT�FӒ�1����!H� ��Y�jI�	3�H���`�Q��A'!\�����:��"%�,a|LϽ����n�G��Q�E�� ])�3'�YHx�dza �J�*�KXf@G��T��y�O��`�	2�]5��,���6Z"^���?�⹀�I�� ���;ϫmy�7����Mgm@�&=��}������P�N1��?��}g���a�KI�B�=G�*{&S��J�%��!8�|�V�����׏��%�G�Y���2�(����6d��3���L�T�ٗ�cʩp^D�B�ƀzY�"t�^��V�-�O�����W���I�ӫ�oI;�~�u"�P8��PL������"h�h�6�o�:����?`�1${"���2��LWH�w���D �Wy��%K�hqA����ȳXg(�@ ���˝.��k=���-��_2��xR�
��4�c5F�j%�ؘ�77ir������F߈�jc��B�GN���f���1�k�+�)��A�� ��&�+��
F���Crk�KR�3(�e�3B#��#|+9�g�d�z*w!�`]�����a�
5 U�k�r2�Y9�r(>�t$�H!j���&�:�"�Wf�镾�*��[�o�ƌ4G!���,���&�P}��ä�z(-���TW�p�������r�����R|?����Baʺ��$c3�s�QS����Z�\S(:�;۴�i~|�LUG��^�Y�� �02"�M ����h>����+�S�<U��������dx��J�	�~�>�.�<�!:��t�X���]+O��}!dFr	ۉ�w����%���d�ʪ����]�xoRj��<C[R2�o�N�#��2�]�������@lw��sӐį.ǄP�xB��;ה��V �h��zgB�� �S���@�Cz.&�qW�K�F��\+����ո)2�Q~�ba(��̅�:�X�N}+T*��s����z���kY`B�b��b���M�����*H�~''�n�vp�A�.���>�q�X��`Ԓ�<��t�#-�XL�B7���2k�rp
��C�Xpj�ˠ=bl��P}r�36i^8�]��P4���Rg�4�1kSJ����|�S���8���#5Ƥ 2`VP��\�#�'^e8$J��� 06�>��גG�VU�@(G�:�kH��S�}�m�c���+��Qѥ��hsf��\9G���'����~�1�)TnT�Mv^������"
��1[ܶ��|�g]Bļ��K^�k�aܺfB��Y3J?G�>�N�I��Oaa�Ϥ�Ivr0;%~aPݍ��qǓ�R�n��OX�cI(/�Nhk������gG��AdRp�+��~�ܪ�~�N2W/%E�F��C������I񧘬J�i���$��ddV&Cr� �쀘T\B�όd"�#�H
�w �}�3���6�sبe8��,imw�HjN��
j� �;�6]E���Ń4X���D��5�����-�sn�쵈�t��Ʈ����� '(�h7w�QÑ�b�H.�j[H��Ygl#ݚ���������A���"ʛ#˼�#$��(O�0M7iX�p���a�e�S͓��qyR*K4��oL�"\�["�-�NG��=��n1�?Xy�����j�Hi��N�	�Ā���R,�LdI�3j=ٸ}�ǝ��:n�Dqttˇ�tc
���T�a��L�tTc4�>�T��ߧ����A�."G�?AR�P4�5�h�P�d�}�~������pQ2�F?�u��G��:� �2FN�V7��WGD�++�^<EU���Zź��g�O��ki�f�ϩ�.Mb�mz#�UoA:D�V�s�E�+�5=�#.m�J$� �Q������m8G͇���������1�������0{�d�V���J
�#E7�̓&۵�q�_9���?3�g�`d5~tX��1�X��$Lv��s��k�-5�um3�(̿�r67-^�Q<?-�+�T�j���\�y�;�@�I��CZ7j���+ȓ0���ӱ�77lf�n>��O����Ƒ���S��*Ͼ ���v�����v����xa����&��5�o����������h|�F�n�����T��7��SU"фy��[�F�����Q�)�ptځ%NKM��\��Y%���Xh�h�]a���<���S���*�&0�eweP��M(����qz7��|0K�0��O�4�F�@ץ̃��f��Ǡ�Ý���n[>:>��V�^�L�1^uUq$�p���?�)_��j��Aq�-�q7{ '�U�oM�b �		�$�2�7ke&�!M��}�M��2�v�w���ɉ��M�޸T�J�rY�q��/QeHP���m����~n4�L�W��E�ac�6?%Ĩ�s�ۮ���Iz��v5ړ�ԣ�4�@H�I�~nd�碪e ��j�������E�9�Ъ�%7��"B �����8��3xK>����r�N	
��I 3:*h�����"N���c���2�`dJWV �	I�%�t������0L=K`<:��Tѷ.�z/}s17#�����<~n=�������ݒv��m��:���ân  dyu˲x�s���B���?Nҧ����vc�i�����7]��F��>�6T-�ё3Z!�*o��A"	wҪUO��V�f������-G�ls;��܎���l/k�`�����aW8ׅW����u�x��|��u<jC�JC��(ݓ�$ƣ����x��&k!�&`��G�9CWg�&M>$eT�\R�c�UhK��b�t2�4m
q�"WtPV�x< �`��A��Њ�L�_t[�n������*cM�mʱ�����~"E#�US��W�[�8ԁ�� �.��;
]s[���V��w'�^%mI�১p����r�춪 �D�
�gwHp������< E���ss�P4�A�+��֯a|��/M�i��,�<�������e������L"���<��7Sl4�gb�/��	�kh�9S����e9�e�&K6��Ezܽ0O4��ph�Z�ht�Ԡ?mYJ� ����aC��K��so��,��
1.��B9{�s�<����Rpm]/г�D����	؋��h���<U:|Io����s��G��K��o����Tg�I�߀τ��)®~[#`�PS"���h��D��L�<��l�ͭ��;aFUHš��7��PZ�1���I�r11�Bq���l0��ѱ
��V���ӱ��K�a:����~!a�6���&��w95hHn�S�6Բl>�a#�%L���e�9�6^|��H�\ߔ�E�W���N�NQ�3���j�yə}PlI@2���O���:V�"H���@�o9��A{�E��~�%"H\B�l�H��^��q��Mv��z2=,o�hT���ELC�bBA�r�d��@^笧fUJ��>�N��������F��Alo���, I=mt�����;�;%_ު ���ʝ��݄��n�������C�ld��������X�������\�ow�b����D^���o�2੖"��8�n�S_��/ׁ�:�-��h�~������a+��$낰2K��r ]�W/d��P<g��Q6�f4,�L�G__���O$�a,1Kʞ�"�]�?�2�=6�:|k�)9��a�S�f�w�Ai���t���.\�ۗ^��k:�j��d,z�s�����~s˒;-�E'��F_׹�XBڜj�mhy��ъ��n�y͢�? �͂2��Ȅ��z���[{��^/<0�������"�j�i��ꆩ���2U�#Q*�Y:�7��oL��"��r�76i夒����b)|���}MR;���ص�P�=v,�E������쉟�����܎RR�I��{yȥDh��:�1#-޷b�2������ I9�X$��\�kgT��ϐ�]� rw�v�T�$#�]C�N���/t#�~��o��r
7NY2p꼶=�f�ݩȕ�eRALP�BkŌ5��*k:�]�[�Q(n0�]�kf�,��I���ED?���<���Ѯo�E)�ښ腴�#z%Ö&B�j�D�� R|om��_c�eGrʒ�����]��d¹t�V�_��5Ψlϒ	�E�������b��D�k�?����@���A���&���ξk�J�ǭn2��a���{���E7Y'U���_�M$9�����h��1�J���Z��1��o�~�m��}�=�L4�U�I�8V����Y�:��Dԟ�^���Xj$_e"J��.��g�*n[���K����:P���~5-��U�j�����R��z��)3Z	��A��`��
J����������m�d��D��R��O |1!i�w n|�Β��<|wƎ�����G�>e�axG]�Z���i/W��@���}.
��?�O�;�N�>_���A_�"[���]���w\��"':�[�������l��^�ȳ��9C�W���}O�jB�����h;yѝ[��l�v̕�M�d�e��%�� >��*�iI���>���ĳ�됉E��0��õk������]��^g��I$p)^�I�s�ߝ�Olq�h�L���L,P�v�ե/��tic
�K��^"�t���4ܗ~"	�0��V��xt��'�)7R~���P�K��fQ�7m���^�&)����O����}g!�}�͝�x�o#  s�w�|�d���.�Y6��,�[ĮH�j��Ս������ ��YF8�..����;R���%H�q~*��R�B�=�.R,��bb:Mr�
�u���9%L�6��_�eoc-�v�z�8�ۚ�8 	�?P��S~�2	/D��V�E�!�U��M���Ts ~P��Ǻ�6��H�`T0����G7\Ԁ��3x�`�8��%vL[�����ڢ��,6vf�i��(�1�j6����g*q[�k��W�s׸܈خ�԰%m c�1�һ�����KIA[?��V�s?ia���\��{�+�����	�v��u�y��������9yAN��DL��a����V�F���7ys��C'\Z�7��h����F���	S�9@��6��1�/�e��u�L�,�KTk�p�ZO��k~�4`ٿBʘ��L�?��B�.�����$���I�z>������'�4�c���v�s#1[�i�{�#�N1V�Dd�.��N-Kd�0 �φVF�O�P#��-�u����S9�^u@���)���x�3�o�A�j���w�+\�l��ѩ'�+X��@_�"ΖY�8⩚,�$��CM�n�ǲ���Ǆt�Atv�08�� �M��:B�s	̤��/�5�R�N�[���7���C?��ݡ#��8\dh�9Y��Afv�7[١_��ÚW3�g�!)p��<mp�˒����T{�G94(�B�x��OK��b� e��C�\���1D�P�(߲�b�?��		v���d��G	�Ӳ�/s ��,N$�]�mR)W�lL�?o���l�G��u'��)�
�6�veݲ�(R�rt�w�-���[����J��"sSi���6�2/���G*/��n�IV����� � �3!�qT�k�kfr&Y�Wkc�Ie(�J��ęυ�����z�0s��j!��Rvm<t���G�	mB�ݧE:�g�e��ַHZ\OuY� Opy)Ȥ<��7���u� �m�ޙ�'�����6M?O�_AK�6���mU�����'^��~jW�Dn)E8WC+Ӗжu4�fZ5�-Te?Q}(�KV*9�S�G�͞Nf�P��ف���_��.�eُ�W: g������(��#.�/t@W?����� ?SE�$�+6vB;Y���Ë�B-Z�ɉ�Ks%�om�h�Xن�'��T��l�ξϫ�����'��,�
S�J��'.n���)m�����FW�	�W��3;C�H�ݙc�*��A?�1be�wQ��m�7P_r��fr�A[�qR�+�5�,)�|������a�b˜���o��9$�g�u�-?�x��E�m��@������m�I:����g�׉�����n�|K����@�?dFh̯3ȹ�j���
�f�юt�P�=8��I�����H����IZs]�:	e��}9�S����ȳPaZ#�[%q�pϥEV��edp'0˄)�W%�)|Ҕho=C;��6���)��<�n��s����u�x])��#�����J�7��xnGDs�tFI-��<�S�����Cٶ�x/�]f����)ݞ�@'��X���ԿCH=��}7�d~���C&#4�LP��[sU"��@}���?�'c��B�#����M�����dr/v�b��/����cM��C� ������bە���0�cd��<�vD]0%�ߤڸ7��m�ݚ��̓9L��˟'պ1L�.�t�����k��p�l�Y'�^�@l��??��apՔ�g�Q�,��a.`w��Od)l.Zd�=
��+ q5���u�<b�������n���%v	��_3�ύ�>S^��H�����A�iDZ5u�`q�0�h��}3�ߓ��CIi��b-�68Z!︾��O��ՇД<JO����䲁�����ȕ��㩚�c�ҏ��e��ك�	�y�`�τ]2�uD@M�y)']�S|y��Q�:�8�
^jX�>�y4l�<i�f�Yg�(sNzʆ[����T\;^ ��֙�ތ:���w+��v?XK��;�^c�;E�/\
h��;������Z��:S���s���<@�����M��h?(��O*Hsc-K[�J�0ү�"��d�?�0]����I�^��F�g��ߍnj��+dҮړâ��)�L�6>T�O��*��93�?�7u٥�X8�}N.���v ��'c�
�f��vX��qhC���E�n��}~����:�JK ����ں@�ז�1}���`��Gޛ3;
>t� ����,H΋{׀)J��g0Uf�^)��i�]�����<Q�+Ja��v�c�I��iw�I�Ɍ�U�VT��bK�GHt��^b�^[_�����/�:1����זu���&����詊�zmZ�)no )�Kb���aXz`ӑ?UG�k�if�w��|�v���h<D�ps2�d3D��"��Ų��!=3o�*)��L� ! A�����z��+�_X%T�L��5�TȮ?떴���CϺ/��{�C��E�n�Au���\�"�^���u���	�b <!p|����Xu3�YZ��vgƾ��jVb�/�a}(�X��J��m�����Ԅ�%s.���h��S� ��/����(l�����ٞE�<-ǩ�ue29��l���5���(�ɳݙ��l��m�q��A�ަǗ�CL4+��	���J���j����^i�D�*�qB��R""FEb1\]�$E�?���iD���*� ����jI��H3�w�(p�V��})�p;G���a�_���@,$.�4����aNCF��KQtC�6�g~9?;�hf�+1h��ĭ��Ҙ"�ZQ���oLk9�ߴ3�����H��,j�@����ؕW�I�X�{=9�m���[l됝�ە�R�C�,�tu=���r;��|@p^�V.P���S9W,,��]gЄ�$%�r�ʒ VG��dDe0�j���=6m�<%2��o�ت���٧t �A.�
�2��E/�E濽�ɶBWH �w�8L0�2'q�9E��Qe�kr�� 
pׂO�2�o��������v���W�ہ��1��}}F�vȥ�#?�S�٧�VO�!8�)8���9��\��B�@��te��/����է}��!/��U�s�3�4��Z�w�9���e�f����$���0�_��qԉI�N`��]b�iXRʈ�
�}3Mzs�a*0�ֶ\0#B1��ڧ���vH����a:�Zw�3�a<��;�uA���")�u�N$)w. �p
���rcA�ƆТTm��Jy"�Rj���־/3��K:�Atx2���\�p�
S$��_E2zD9�T��FH���C.Go�)�o���h��I��q1LHHV���)��!��jGO �y�x8<H��M��E��q:�uP��f6�����.e�Fs?�!o�a!&��M@ ����N,�~Oߧ�f�8�<��r�Sj�ļ�S���qm��,�΄�̄��,���O�{�;����a&���I���t�fo��b�cV򲷹��z��/�����ڒK�w����S4�4���{0�o�ʢ�z@c�*9�=��q.\ܹ�}4�sI�j�h>)�ǟ
�1����3��<A�Һa��uw{_��w�V���𳉍^��^2m�����I��P)���z>��,��C�NŗbƝ4f�:٥ٿ;Vkn5ނ�]/�6�h�z���-y@��0�?�*y�T����: ��2�9�k��ڨ`�_��{�����~~զ!�M��^���j�fO�Y�Քb�^6<���� ��<��P�jb#��,=���]�L,��70�en�8�t2Ϳ�1Q]����Q�+>�a�"Y��f��	�c�?7;E���0�*��'�W-բ���U�}��+�r��b �d��SH��u�L���e֢��[ �BB[g
�����v\a�7ht�Ҏ��f��o��fv0.���ؐ� +����َ���C��|�a���O������ ��@
uX�'_j���w�YN�w�
���3�[���/����t�^���j�xǂ�\��m��RVc��۾̝���8�	�@>)'UU�6B�IifJ��X"�����!Φ�b�Ӑ����^V9�nf���V^6��Y@1�@'�E��u��d@7e86 V^o/��Wgm9�h6�db��*(�buY�ۍ��r�uJ/��CD�W�^-�N��N�~�Gf^�G��RH:�g��.?z�͈��c��Wυ��^�c!� }���7I�N�6���9<j��6X�8У�=v���?��x�Ĝ� �/p�~���AѨ����a��Fk>��PT���G��4�q����~^�Q���q�{�ɚ�g��.ҋݮ���P�U#j�m[T�nG�!Qj#�>-��ҽ��ÙwfYF���H�MltO3q"��;U5��uL�
n[���t7����j(Ng��׼�ȧF��j�kT�'X3C/]�޽�\sd�/+�7�ve�t;#`��JQD?��Z9�1��������N{��w�(��:�栨�B�)a4X	c����ř��7�q$�ӏ�x�|D.���ː�����fqh��E���@tBF#����&�$2��갦k���-����Ѝ"ӕ7�������"OD�aM����{�ZФ�u*��MᇟOa:T7Zx~wI=>��gS�53��PMIUK*X�-���D��4Dݚ��4���7�F�ܵR��|���.s�΃	��N]�(������j'���d�7�R��H[�Zi��r��8�9LW�w��Њ�|r����@A��p|Y(q{��/fK�)��tݢ읷W��ҝy�օ���Wp˅M}�7��T%B^'�i^3�,M����G6��c>�J��ձz���LiT� >��А̏n%����Up��A��ip&��v���w+v�!��X��a'X9H�&�����S~\�q�fO�FfY�L�kM�$Chx����7SZ�n����yX���I̲�L���='6x�UIk�E�4���l:R�%���#P��=q�5,�Xh�[�BBB��1A4i�;�g��X�f���»��z\�����u�`\��� |__������,R���7����ӪK������:��+�������[o,�#�y1Ry<�sDb��9�WDQ�t��$Z�x/���pO^�0k^g����o��K�%&��^ȒL
V�k��c釄<@oM�����Y�2:�Q���r�����Xܞ3Vȝ�z��R~�'��	ۛ˗"*��0����\���{�lMx�]M.4��b���3�)��Q�R��� �&�Ӗ���An/pՙ9$��mq�d�S��?��a@��6τ}R�z�w���]�Ҫ�R���LlSQ=#�� ӻl+���M��*�3��ƪ��k�
��g�M�P̎���ؾ!1�Zhܑ����#���&�)Sۆ�Cc�����<��۠S챩����B�S0$�;�?��q��r3�A�TX�q��ȕ"_�Z�sΞ�%��P� q���od�:�{B)q�]�Hݞ̨F8�*MظV�#"����=V��`�&g���{� lK�J��pK��Q8E-�c�h7��RP"~"��I9.S��4w���%^�Ỹ9� d������'���p�	��:�{V��`�!�צ�0�T[�}�� ��g4 Fp"ؾ�^Ac�滹( `�d��9j-���t0��|�f�{ۚ�tL�E��"+6�g��d��4����Y���f%��Y��.wu�:t�O�{)&#g�5�N$���($��i�@�QFƛ7Q.���\�b�'��26�W�&D h�K���!�l8���G�)�G�� ^�f���ozKc*��^��]9�Q��,*5k�2���i�D�￫����U��Ѹݍ3��z���'P���"{�J5Ē�בL�J=��)n��d���e2v�fu�#��w�G�5�z�@��R�W˷Z�2D�F��?����8�k��@�)⽬� �,�񯸠��vL׻]I�y�O7��-���DU	��*�� ^�4Մ:ZjZN����zU'���I�XM$�C���Xk!c�jݦIV�R�nO]-#L�R}�=K�o=e0���fw�y��ԦM5fWc��Ȯ~�.��*�3��x�؏�y��A1� I1��jd��i.x;ze=�P��2�d]��z��?j����<.Zp�N�H50|�D}c8qR�k��j�ݴ"{ݼ�3���YF����\��>1]�Kx$��.`�ÿ>����u%b��Ī�o�>��%M�0���������*'��;@��o�S��׏E�dQ� ܌�5��>�&�ĵ% ʚ8Y̓�7�b����h���0mC�M0�:��Pv�����P�����'�m��NJFC�pE��zU�l��.~C���p�$�̂��ч�`{M��������8<1
7��h�l;c�jc�*�����X��3i�� +�ø������y(���� �[�cȅ�t���@���;�<�l劕�_/����
Dfe�AX%�W+`o�wF(�&�ΠoǶT���5	�P'S�6�&֘|Yz�L�?����sC�U@��e��E��OA�2�w�|���)��W��ݶ$S:%w�,��PlO�H��Ld���6	\�4ò�q�F�@y>�k˫)��;��2Z��e�THr�(8�DU#�G?'e d�@�w6�A�A���ھ���NLІ���p�N襜��M���`K4Gal��z ������tH~r��(m�S*"@M9s��?�M�L�3a�o�
�����p�����j�^(�p6
�2�+��̌Yi��h+�g�5C�a�t�ZoQ�����̓�be�?�9���]fp�g��ծŁ���┳�r�(:��r<5=����^�"��'W�r�1���\�[�9�<�D�6��YW{ၷ�5����H}7Q�VK�����E:��f{�HS�f�����W�׹X��f�!�]4r��W'ΝLaf� K@�	��OޱذN��b��,oĻߊ�Y�.rAV
�͒�x��ߒ51y�2�?�~�����lW�����;ΓMTR&��d$5�W�����ε�b0	e������l�i�<���^.3Ȧf4��02�E˵�I�lP�	�6��6�Q���돲,_����޿W|x��~�2.�׿`TXUً��G.<���� �j����c�I�]8��
\�]s��Z����9{o)�J�w��z�攺��xe䚨R��Ο���7>P�h���+�N�"��"�:hI�����ŮF�����B"v��3�2����J�IT`ҫ7�]3���/n�bE�98������rB�������6��봭�#��gBF�F��L�P!��
�=�7��S�X�}�j
���M��GN���,U6�b�o�{G��ս.��TAo���H��Wˈ�$	�ϭac�� O�t
Ā*j�$���z�*n�t�߽?�r7��v���_[��Kf���
[2�Af�m�N��m	|�i�\3q&tY�ԩ���k�:�R%�)�%�
�c�}�Y�=����p�`Es��/�3�7�ڒ኿�2|Z;�yk�$����V�>��}����7����tGv��~�(�Ke�h1������K�G��A"M�G�/�t��y�}L�]p���zf���>��A���jF�3`�G]6��pA�(+?�b�O�W�I���?��|��R+�<Ɲ�0S�7�0lF9���!��+pa�yН6��M���%J�L{6$o���X,^�'�c���D�: �A��}?��i)�㔬)��D�Y-�r��!�;(�wt���D#ͧة1�������"���-��H�0�j������)Ц��{GǈS��l:;�I�s\�G�'�9oZ�K��x�]�jU&�fj�M���,�'vP��"h#wy�2�:M�������,-����!�K8��9\�uD1Sߵ�n���L}jQ�^�0"h��~��po��]]�{u�6G(_��P�h�l��"����:�]��|�W��Y>*qѷ{��q�q�$, ���{{�0�x��c�P[|�x��0Se9rα7C�щiq1�t}��4��g�qȼ��
�W%�lx��b�2v���{��v��\,�� ۚ�}��������V�ġ�1���_'��ȏaf��WKG���R�@�RH�w�\Ov�'�}����G��D����>�E+"/B�@��0�'
JU�T��Ip�\7T�N�6��k��61U�֧�5���Z�
n}}B����t��Q�䤇`�+�@���+0|�%��֩3�kׂ%7xn �!vO��T�?s|��e����+
���f���؄�F\�O����ͯA���@�a�	�O+h��ծ\F�. �ం�n�?E7�gRa���22I&�e*)�q:a��WQXY�?��c�T+���x��	>��`�I�du�l���1���f�m�A���6��)���H���	MR^��4j���F��\�`�R=.���6{�H_�͉���a8"���B@�Q�:k����(�o2沢�i�H�l�O�y�w�q�a𝃛�a����wc��BHT�H�(�Mbٔc�fw�A�0�t#�%�]1)8 o&���&����z��Q�;@^7�
&����d'�?;����A��o}���μ���pT�X(�up��u��~���8�ޖ�+k���+�o�9�'!O��\�o���fH�֙T�'!�������֕D֥�4��_���/��]=x����E%�3�����p`⪚�I��>γ����w�~N�?�H]�:(���t��	�$�?�{h���f���J�Ħ!�y����=W?ې1��W�q �ۺg*�ySq����)c�za���Ӧ,�_�Z�C���+�a�ٍ~>���.�1՜�X[`QIST��9En�Ƴv��ޭ�k&y�9��#��:�;��%LGLȪܓDY���z`R�/Rs膢m{0��+���T�~sd�\�ڪ�|�4}B�48a0���62����q!a�6�-��v��$�����E�`�'Û��$'x���Q�5�а�=��$n�N<�$F��z5\$�wb9�8>�!|��E��y�U���F@��7�جۙ�������#��F����	��� e��#���a��<�3!���)��S�
-�tSRX��K�����D�ŏ��D ���wT+OKKe���+qk�ˤ@qOu�4첞�ήBd]W�k��ƐJ�SGNS�� �τ��)�}hٍ�@3��>8p��Rd�yk&?s�ꁧU �h#�T��C��A�O�E_�;����M,p��AR�[� J:��L?��6^]��nѶK-5!��S��a�_+l�׀��(|���6><�e}C�H�&��^��[�+�ӝR9�\�
���4�*�Q�
c@(�!�k�͊ݪEj��U�K��L6��C�h�_{V�E��Vfg$s�[�o�P��o�+ �q����L5~T�U��6z1_5y���,f���HY:��;�1:~-dX0������``�4¶�k×�����O׋5iB�.s��2+��۽n����<���$4g/����t8���Ŭ��B�,ɷG+��X��>�+�꬘R�i�D� ���,ʶnC������u*T��#�����]�A�U(O�? �ׄ�@C[��	vs��IK������j�^<Y7&�h�{
���c"�H���_3e�hUHS�;��[����4g3)�=Fnk���������[��D�"�?Lӱl��}�d�8�!��\"՜�Ȩ��]y�\k]����"S�dN��V,y��=�S�♹���C�U�m��.��;��3�Fv��������u�fʢ{�>ʫ�@��Ҩ�z��!l����ԇ��T�qv[���BS{�V�Eʿ!利p�t�ؔ�`��A,������qE�Ƈ�^�U��YT=��M�8O��b�6�i^�.&P� �p���܄fm���-U�p����`0�[��c���?`�f�˿�֔]����Zw1���^B���v�W����9�%Dm�7�>5�87�4|�/��#:3=����V�%��kM��_0�b�M�a����w��96s����9�%��!�!�v�pd���j�Y�H������_�O����-��0�4lw�����$|��YL����_ܹ�Λ���"�M.i���LE�L�/Sxk�Dc�J��֘��!��|{ʭ^q���P�r�h���!fTTu��5|��k��\ֻ��R�B����Ӧ�	�����S�3EOe�"��E�f(��3"vg�t��Z� ��~��W'sB�t&�G��q�r��{�S迱q(�~,{I~�r*D-����E���ÃE�Rq7����bҁ�e����h��Y=5���6`J5arH~���ýik��(D�i����S��+���[�W�]��y3h�̪a^nt������M�1�@�"�����|	�,o<��ሞkؿ��9Jĭ��� ��o	��y��^�JRg���So�쏶r����G|{��WX���N���=\[�k��xXJF瘷yP)(.��h������g��\}�Z ܘ^v��S�p���p��e��)� ��j���U�@��~�raR�T����:��=�����/�º��C�;EgM}��K��^b�֥���qc�-�xY���hu��2m.��TyN�P�c�*��*���
Сr�G%LD��Um[Zmy�m�����ڪ�v�bc�H�5/H.~���..ig�b���
5�.y�_Ւ�@G����Ԗ�)e�V�����[��x��g���=ـذFM��ܬE.q#o6Z�iA-&v��cG��������d>�e��I<�W���ɢARB�彮�cm"�VLS����+^?� O,fr���fs���l�}@N���[:*��u����y�9�g�у���-�vh��E�',�/h�x�b"���ڿ&M▫��K���,O�����(%�g�(���8������K`�b��ҫ��R�gȜ�W�)�b�,>���O���⸏��@��}��(iF2�������֮��њ�5p���e�����IP���������aAU`�2��ɞ�	%�_�o�1��N伯SD�X��I��9(�q�8�ί]9A��}�Ё��e���oAB!� ���ro�H�-�ÒC��o�6J���3� ��߿��ޛ��:�d�XR%B��N������Z���A_n�V,�v?=�1qz:@O=�R��E���<�z��>���f힪������$���R0�9�=I�S>J@U��o�Wv$����������q�|m����-9sk�����pn�/[Ϋ�\R�vC�M��ж��S�r�1p����̤�iƷ;�E�+~�K�'��*����ɤ^�0!~0x��L�B"AA�-B�Hͧ��S�S���U>���#�����?'?��1�8���ju�,�C�����1�k��R�j������s�'5��(S� ��w�^����R�+��G�)�GH%!)�7̄%�� �������G	-[�8B���p��k��D�xo��(AW�@
��e���gP�¹�l�$<H~���˻16�20dpdS�U�\��៎Ep��[������҄uy���%mJ�bX��`��&�A���6��%ې_�m���'�h�o'�
��<+^�~��h\X��;�)�����q񘔠 ��=�bRYI(v�KܜC�Y�}geR{ �I�=���I�@���i�9���yb/]!�LL��C���R�!Xl4�pn���Ţ��A�ķJB�H-Y��iiemWp�eЂ1���Aq���f������0ه��E7W�J��	O@��[͜+�k��[RE5i�g�z��k�X�ޥ����m�g��ߣP0��	<Y��d� �җ�d"?��ЪW�0�����ņ�	���	W���ǉXS�=�3�բ芜��s�|�me�Jlv3(���F������:%qy��
�f)�`.hH#*�ढ�O�f�u\�DoA�D�Y�){h�,!ޠ,�D��yKT�mz'��<���#�i��j9�b"ܛ��Yza �:��4}��vj��틁;B���B!&tUW����������?�����?��*���~:°��� ���&~�K�ľ#%i���5���S��#��fq��-m r��#�f�H]��೟�f�B��c�.�q~Em֋���;�� ��(����{�ʀ['0)Wj�]�4{�N���Ϳ��p�.ZqY~ڃ���w����)�v-�<g~��8�N�7/��n��>�hN�cLL�p�͖=ȨX�r$6X��{�l*J��T�@���t���'z:G�I�� T��M�.{��s��~�N���:m��,�ɓ�
�Swܡ�Q���4�*�)|ג��v�ۑ~:M��r�$��٨�+QYS�_�GwUk_j/2ȋ*r"T'(�K'���� ~�fV~��4�kwx�R�'�mM������R�����&U��]G��ݸp���r�-q��P�%�߂�\Q�w�im�M�
���s=�$�Fٷ�[�%) �uX�u����W��Y�fD�ǚ��0MW�Ǻ{}@�F�ē�4���MI���~3��9�o8y[~A3R+�>0H�r�L<�e�9�EV�Ϡ����`8��(��E��z�Yt��!�aK#Ϋ�ܮ�Rm�J{�;��a���A��=�@��A�X8�q�dt#��&�z_:�҂�eq.��/h@�!T_S7�i���h�t�\�X�6��	uw.���P����h(��"M
w�ȅ�5�K@]�.;p�TC ����0m'%d�f�N��U@�;���]hj�I�t���b�t"��"}�
���8o���O*>�7�� Qr	 r�uC���l����"��\*}4��q��u�!�������iO�a�g��<�$VK����:
�����#�%H��Lᮬ�u�0L��y���'���_�1�r	�V��7V�]�:K�,��j�R��������Ҳ?�s��Q�������0�����׸Ra 퇛����E��`s/[��|i�d��t(�i�4�US���gd�����!sjS�k?\���(�:�}f����T�!��B����+�$�>T��{�����D�H��g�oi�m�U���{��]��Kk���{б�l7��L�6����$�8�l� L3Os���0��@�b�]!aZ�6��_�9��w>�
$��^���u���y~��6��1�,�׹�SYF��1�~TY�L?��;;��P���9��2s��1� lH�|tL��fs���g!mD�gi�CuegjX��v�k�j�7y�$cI6�qO���ӟ�����d^m�ł��A�b�]P��Y�mRO^|0函'�q�o�yOt�w�[Ū�f��9��d����b;���=YyhFku��ֽ�R�#��Z�r�a���L����9�7W�̩8���Hl.-�k�Y�k6�M���n��!BL�/�I�[��Y����a�S�H�G˧�gX�"z��'f��:����)��ໜW5�@Rn�*���p�-����\]����U*�X�<�Db��x���Cm�$a�EQ�vԩj*�<��CʌC�E�mT� ��Fe"^�R":��E��.�f"y���� ��=��������<�`#3���%������1x�d/��-?�#��,"�y_L��"�7'�w͝^��Ak�|�F�Y��1��B?Q��L�<�M4�IQ�4!��~^�u}�8����ɕ�0N��Sy�mD/Y��s��X}�(}\�Rw}A>I�#���!�y��\�DM�ѽ��$�l�e�t�r�Ï�nQ���#�=��o�����K:�id�]N.±�u�������M���*��h��>���QL\���7��Cz�(��fU�Z��P󫏢̦xkkt���`� GΆ���Y��@�9xl���MC}m���F��x=�׺xX�UL��S��kp|��p���
��>j�T璽�pJ~.����)i)������y˜��̌���-=b�?�S]��V��5�b���?Q��Α�Q�����8;��Xl�"�z�\�Fq_tAW���%���TM�A-�캝���Q*�f?1�J*���?�Y���b����v�+s0�Ee�\65U��ܭ���4�I��f�N{F�*~�w�V�f�4�-#��j��8�yV�]���ÕoÁp4;*�� G>��:�EH'��֤e��݄q��+�8K�+���NrJQ��������������hQ6}�Ρ�D��Ah�`��JE������L����l�Vd��)�
�� 2wUM{�#��|)�U��ϑ���[?~kx+�e���� P
t��J"�n9�ޮ�{K��]$��DX|�k�LPM~�g2sc#o�|���FJQ��P�N�2"7��ke�<�u��F��K�j�M4	ɳ~�L��ǈ�!�OBJ�!k֨U��'��l9��=�������¼��)���x�K!���Y^B��p!f��=����tp�9�(v�j�^w�*���V0�T�q����'�}D-S7�@[f���"pGl
���|ўw�౯�{��W S�ԝZN�1�ŗ(�>!�=M�_Y�;�!20�^���$��h�dw����	�-8���fF��hr���+�q��GF��^�%��a�`a5�0J LCr�O���a�t	�%�]:�#g�vl&6�o�bQ޷�' H�jr�	@�~�N��̡[�mޟ���&m%��q�;���.�N?<]C�� ����ܧ��f��EZ<Ͳ�,X�M[�6�}����R����`�G�T7蒰�uK�ag��t5�T�9�^P/�����bL� ���="�����V���P�
�Y��?�ّ�V���X�S��
��˟d�R� �0ZI<�p%�Ф̝#p�3�J_�d�|<y֧��^��	��3�!BI����b����;��ƣ�5FX���M�:!����˙W/q�;����Y�i��g/�r<b���d+=y�0fc��Y��F��p���1P�aa���o֊a��P��-d{jW}~��1�r%l[$ߓ>=�1��#bU� �ɪ6'<�3ʡ���)�4��P�r��l��s�@���+�8�9�x�ڹr������7m��K�
-�R���U�q����e%�Æ����>h�؎L��a�k59��y��0��Lh>��۩E-�$J;���uB��q5�n�B�,�8�r�n�b����pևP�q~.�!,6�-�}���y��$�%ڏ�E�����s�o�����>�3(e��.��d�P��_�����p
[�ޕ�6�К>������3��Ï}}b�k��K��g�ք\[4U����|���^Υ{���l���m<ZU|LW�/!�+���
��Ѡ�� A���|�4���;z
 H��ټ��y>d��gʋ́R23,�:�AN�EB��yNa���Q�O�hࡤ�n>�@p�O[=��\��V��;/��wP�;�Itx�E�[��+��C�X�^X�Ƒ�����,����TĚ��=����M;=�����/�����Ν�ڙ�Qп�b%H�XO�m����9��	�.�
є�jq��qDµ��K;�1����J?��.�
�  ��(��-V�p��!�oWÊ���cջ�Gli�#����[����;��-�Մ.���r�7�ih~�2w�ۇ�Yl��,�2e�g�� G�;?�G=�T�V�8����n"Fx���v8T�AՃ��@�}�U���=#ؙ�Ϲ�Z.�f�]��G�"�<�Ue��@�6mJ�Ô3�4��Z�b�F��<�B��2�2p#I�x��x}���{�B�>{�wJk6��aN��#gôV:q0��.\��܊?]uE�$;qCC�<#!�N��h��Q��V�Qf1l��I��v^
m����n��Qq<�l-r�݋������'P8���p�Tg�7��!��?��Z��41<2���y���,'*���^�H�=@1�L󯣼5b�{dI��|I����w�5���H�J�DG A�Ϸ�ZW+s�h-��*,!_ZTzyf���㡶�>��!�l,&�0|]�?�F`�$q��;��	NP�J��bS�*r��S��$\��%5�I7��4@U�N��\��<]B×D�N.�����!��9�!k���ˊ����E_��ݝ�J^ejJ�zJ@��tq %�U@X<D1���Y�s����B�q/g�C�ڲ�ϡߡ�ZdҘ���E�YT�s��9����4�?��rn�G_�6I�\ύ���pg5��ߺ��׿�8Z0��lZEh�EDf�c4IP&����-h"O��Lt,����⾂b�Q� ��]�޳��^tƊa��?�1��+��]�_	��9Q�0��avwɓe��� ��߇�G�a�F�e;:�234��O|������O���b����(�EoL���%V�9%WI�y/U�ܙ��}Sc��_�
v��V�s�S/�l���cW�����j��	�T��
uy1v���R-{�A��C+�%���Ht�^�v͈�`�&�:�[�b�:����w���B�zj|r��9�`��0U`��0a�?�ª��(PL�^�,�Y+�ʠ�%�0NE��'��|N�,��j����>r�W��˵��a��:�>��1|D{�j����-�Y�h�JB��O�;?�Բ]��n���ybU.DV@9��`����J��qLL�;	�
Z�C���ĸXߣ�h��%��o������^7�$��U��&�3.F�j�i��'�i���i5#�Y%j�"��A����]*�g��c��J��Z���(�Ja�j�k�	Ȍ]o�:�]��c���7�(�JpMb~���?����Ӂ_r�?`���8��j��I$�Q��fy��cI��'J%a-x��� 	�Z��'ӿo2��%KW-u���X"T.�l��65bE�5�2�����vB����h���E��I5g����dR*e �`��M���O ��peUh��7U����e�y�j�H�s#�����.�k/�
��?&@
2��(����&Eojl����~�ч�QP��j�����Y��gK,P�
�
���Z��Tb��H���|"G-3P��1�&E16��=��cL�ݑ��:<'i�3�S9Xtu�e�H�����k�_��H�:T�g��dO.y�A�Jj��P��Ŏ�6�kP-��?f�8�1XP����@��4�~;�&s1��bu��t`�+zGI�5�|���O�)kr%��J��)��T�Ʃ�g��k�K�/��$�P�7��a3�+g�+��W���ltx��Z�~�N���FƐ���Y�ԛ�����ܸ���(�Ūu�V@z,�x2Ot��4p�����cp�7�t�������pb�f�w� Yd�p^�G0��I��r�L�����5���v#p���]��KS#y5�eXT�:)6�	0�c0��Ὑ0* w3*2�[^n,L�m�4*L�q�g�S�i�w�|$���G��]���
���L��W�zٚ�	�J2���mO���&Zg���n�d^�����Fƚ�Ρ.�����V�����*p4_%`��@�Y�^�g7|;���w��F��xx�㖛C+�!�+�����+��z�]�f�L� r���B	0�:�vų�J�`#z��<�k�,2O$]ԁ�K�~o7X#H��am5}�W��Jz��O���4W3�+�y����Vm�E��|�.�TQ|%�u��O�Ћ~����������o&��29`�YSj��	XMq�:`���+����dL��������T�l�.E�;SڭqF����dB��D*j�h)��iMm �L�#����Y�Z*� n��vm��Mϱ�tG���)�����,V��޸r7�P�76�c]�k�ş�׃M��	ԁ<i����"r�<�c��	�9�K6s��|a�t�<�ܹk���� �nx��b��x6��m�Z~�:l,���9QU*�������<��a��tM"(����1�A� ��>�
�[#�}��Y�P�E#?>
��Ҹ��%�J6)����@�WH����_���Q��}~�o8���!����0Ϙ��'���QF�֢�xY����$0&�~5�Ƌi�kB����[θ͉+P��wu�k��X�I�e�⨭�F�] U]b�Gӆ���%�J-y�E�����"�缻��>��������]��r���$t)<톝���C0���Hcz�{�R�
��pN��.K	���7щT�>���y0l�d�hɡ*7�a|r|X���Gx��А�Wi��� Pa�k b<~LN�EJEI�~Ԏj�Q�sa�a��ܻ0��{��!���Oy���!��ӊ����U�/^#׋G�7��H��HM�6�Rv�Źg���9q[c�h7�*����nL[�և�V��T@��V�4�"����Q%���Ep�~��9�a}c�{�����L���O��J�m��۫��H�5�-4��.pP���Xz����'�H]xжel��]��މ,,m�e^c�Bӫ�#�9e}�*�)�#"�x�¦'Ti0������T�j��îq���(����e�xt*�)%>C�v۷s��&��Jv����-�0�h����ǘJ9�U\�0��Dr &i�S�|�p�WVF5�[��й!��\?�ƈ-㆕*�B�1ƀ~$X�~d�$��<�C��-������s���G���o���c���3�?���h��Q�"��Q���]�&�F�Y��|5I��lj(]�o��u	x3[���Z$tP:��!����o��Q��u��T��Z,�DU۠��.�d��ԦE{i�b��c�?b'�\�yX���T�EX����h+5)1��Ih���3#c3�뜺�~>-8.�J�����:J�;a�8����N���q:qK���^��wU��K��]���s��ӣjOmob�.5̵��F�9�u�m�&t���(��E�0�e}/�\aDM0OsB����\��(����׉��\�7�KHz�>�*�o*�!�����Os��8�nxJ\z@l��tQ��O�� @a�dQD(��u�9{h��$�����ǀ�xY���ޚ�.Q�:9a��n��J|����Pb���E��M��D&���-t+~�%�izth\&�� ����5�ӵ�a2V�h���qK������fb�3�qT<�V�A��3�ur����Ʊ=��=��߁w�&Y*4���J�e�$��m<B̽�%Be�#�#ת�r���s�%K�\�Q�T������Cm��a�H3�����H�<y)�����	L[1%��k��
z�=��L���thC��H�0u6��h��Q
5F␫�%��zO��Z���.e&�O �9-\�sBG
ޕ��Q�6]ƹs.��uC�=�و?�]i�5'��!�Ya���D:��nG	�9�@����F�ɗ�m
�;E�g�� ���i���Up��^����j��0��9W���^]e��i[H!_'� �?d�}��c�;4�O/(�-U^���E�w4�P�|�p��
4�@˾%�e��>��~���w�q��«���A�{��z�u����kǥ����oH�h0ƨ�K$��2����7����_D�C�u\�w�������=��9��I���N��pv�=Է�`R;n���:r=q�
A�;0��4ϧ��,WI �h^F��KmD|��>�Y T��jtGC�I!�}��8��92�S��������aeWػi'H�Ni!�� �V���] �#�<����8D�wCd��M$7��	��T0ǹ�����s-ř�����
B߷��E����+7w� �v�a/��������/Rk�
$��@-�9Q�X�7*7*���ve�y��fO�4���s�`�8����ו*�8�|�����/C��82��<���-�#�B�����o�E�C[�܇P�z��xS痛kK�%ݥ�����T/�{ b��B�߉j
��̰+r�jYY�����_�F3�o�<_��R�:g���_M���j�N��p\��)h^�d\<	��Ƣ����y�euȭ���	��^�ɣ����d�&�6�Uo�����Q����0��j`�W���\�O@>#��y�ǉg�x.������ޞ>2p?&ҕ�/�ʙaoq�~{��&1�C�mǢ}ƨ+o����:�K˘��J:�C�w��"�XaV���er�qȌ`{�4�*�,H�5��}6�ćf3���x`'�+{X�ϭ�DT<�G�^���'4��;� H�\����5ʚ�u�$��.x�>��:{C���->J����KX0]_��e�xƾ�Ne��ZG�3kpO�p��"�I�A)��A��S�:Sqa��mC��1\��l��y����:�K��z)�6�V�!E_���Ņ_��hPۊ�0)1L�=�|Wv� "�#yJ@��ȞKȄ���a"^|P�s�^<K'$�v���S>����c�@|��hAH���ojͫQ�����T����_�������L5^^�ҹ>%٫�T6�҉h�w8���"�5�r��t��ѻO�0���l��Ԙ� �;���I�� �([9W.�Ӑ�̼���1iU_ǲ(r�X����n_���^�Z��`~��v!�Q-QG����E�� dUs7��I��V��N҄O�q��,�?�KF�%$y���C��5������Wͩ��p��AXM���}�a��nNH�q�Xb�ߤ^������ ����IA�p1��á�_�%���> A+�߶��9���N�cZ^�P�������\�NM��:Q��\�	Y�<�$�Y�������������۰'�	��Z/)'�)��ag(�y�g�N\É��O)(��Vs	e��m�J۝���!��LDo�X/�$‶ۀ���
xN[t�w�z�vݢv*F�؛�i�D�F��
x��%I�E�+s��b������>���\��yrBV��?yyS4$�D[J��5�D<g�잟r�UE��Y��ۊ'��W��G�vd����7��>��6� DF��?%E���y��ʾ��{���u��;0G�l�bzka<N3�����!ni�(�5[>�]%#E��߳n�|t�����+e,����0�c��Cd2�{>�{V�{zѐt�^�ik:��h@L��?u�(R��/�4wo�p��ߦ7��y'����h�
��,q��&�z,�U��߼�%I���2�^ [^S	���4Y�{C�K�\uo��H��3�+-��iS�V��
)	����f�o*�x~�Q�_��Q��<�%�٠Z!by׆E�q�/0d��N�ܝ��*����4H����Y9��N;��Ў�ɂ�v9�pB�����E
 L(�ke�|d|�k�(Rٚ9��M�m�C�Y�S�Ja�ќϟ�$_�Hb�.z����%u<�% �=(�^`����Uų��&��\¾<O&s!��2zy�kp{~�4��N<#����6�����G%�R�N8Yzn1WJ�����F�R;{ȗ�z�!���s�F#X�����YT���מ>Ж����������i)7��&��ndϯl�T�Ɛ�o�C)�3�k��l�s�9�.�'�����k��o[��N$�O�d^f|��/��AS<�Ѥy���`����ƃoMluB��C�js�+�
+)|x%8��lU�9н�W?��-��~���T/\[k<�郯l
ʿ��aL?[�3z7���<���,D����J՘l�a�T�}/S�P����̈��	�EM��U�ߑA��b_C.␘�s��ް�)�12{3br8�E�������'H�l<��sֹ�.60�� �?[������kS�Ac��4��M�r��Mك>P��$7N��4��e 'NSپ�,�>���S �՞h`�tk��bR#2e�@I�oT�ڭi�QK���jۀb3����x�s��s@��p�օSP;Xq�|�g@a��@���I)9N/3�O���.��G�@�A ����VD8�V��Ջ�L�'Ѷ@xp8/�X;�9�� �`HH�eb~O��?���t�"��p�[*�坾r 9 �G�.��!�DzɚI<�>~ܶ'A�$��vs�K�<��=X���I�LG��C-�p�O{c�o
~3a59ǹ���q��q��K��CX2ؐ�}�q�{�P3�e�w����["�`�\�_���� �3���a���筎���6e뇫���(EES��P�NG^2`;�A+4����6�z҄����D�w�F�j��'�=Q��Ii�K���?���v|���Yq�Fop����1�ޫs+/��l>6�#��_�g�mϞc�=T2�`�7�K��S>�Z3�����(��D=����&^E�6�":K����B0���$�s]tYsT=*��š��!p~2�Hx�d�gmh�H�m�E�/G�� DzB�Щa��O�JWa���A�N��ʳ�D`}<�����]����<�b=�;dG��/�сwN�ݗ�'ʜ�_�?o�W���a�7hmKvF^MJ� �H��v<�����I�~(RJ�
�'��![�0�<IeoJ]��S�I�ꓢ�[mx�vn��P����@Ea77ɀ�l��Z�y�O b*&�@𬃜T�UL����,Ua�Ne�~��  �ݬvQ^�����_�� ל��"��őG0AS�{]��v~kTiux��F³<�8��}Y`�[�緑����T�~;;5�Dzr>���8aw��bmV���
Vd+H��mmʃ�+�<(�]ĸ�Ƀ}�!x�ZĈ?G̡$,P���"�W�),Azp�e��-������*�E�_�^q�^잦?-���mh��0[��"XYQ�+i��+ܭ���{�p��~¿����H�d}��oI��C��8�ܙPdJ�,�� �u��  �O6��7���,6�U���1����Y�	��D�0HM���T��v�)�Q�cC��=F��i��E�NSL�t��M㢮8�b�:��w��)�97T��*jf�F������������X�?t8I�8�%覰�=c�-9��>p���56�[��׭�mS竿	���1��9l�81��x��9�-v��%P��5t�=��?{I�����)�!��T�kį����P~)�������hOt�dd�p�w�cmK�L��:Pta�RXP���)(��H:Q��s�������3���)x������AFl��@��j��Q�Q�t�>~ъ`�jfP���:�&�@�h�#��7�C����9�;��Wi�#Vv�������}]\a`a�P�k����:��r~!��J����+�����4o�E�5j���Vė���gv��}��Գ��lƌQ����mJj���i:5�S��h56]���������\�X�|,R�_F�oxh��,�@��@�wn�I��g����Lj��pU�؛����T���,�Ͱ�<�5��w��T�w�D��[uQ�|����Y_�N))[酓��{)�N��"n'�P���M{�̰���#�E�Ǵ���6�>���8'j B�!�e��$��L��/����<�I@�~��p+R���虅^�� ��;�]C_!c ��%�s�.TYuR#����`����n��4�X�HISc���_��i0h㗮�
����(�����"�F�w�n�
��o���g�K�,��(Kc��m@K�׹ �׋c��I�j���GT���b�*�\�1e�
��e>)^�X~w�+�4��{�Y�U�Ċ��x�DD�A�7V4@x��� ��^Q
=~x�����]�hqΨ$�A��ik_����k�W��hS�AF�a��؂t)�� ��	��	2O�9b��(AIt����0�C��k��\,3�b�gpDqh{ٖܶ�~��L؞�Ce��	��ꟛ�c�k �!
e��m߫����aq*6���0��F�7FE�}�i��޶�d��ׅh.�DS����C�Ll7M�t�~�͆�m���M�3,/��糡�(�? �L}%�%�&8D{���bܽW���7��R���<����g�YZ	��õ�ށV��'��u,6����������x8�K��EU?����|��=qX�;}?!��^mDr܍:hؚ���{���T�+KSLJQ�Ý�q:Q��Vm]��n��s3-x�Cl�'ʰf W����������d�(���M�w���e%TZى����9P�hT�A�+(��l���E_�t��I����9���]0�60v�6ۻ(/�pK�o�;�uN�}���O8�^u*�wM��#� �y\����C�>��UK��$�t�^����'����>����]`�˄���zؖ���6�g9+�"���$�	�+�}�6��Sa�������Ԣ�^�� ��^��E� ��Hb�5���e�X�ð����Ј<(7���@�L�Î��KО��P��g��i�#�@��g6Ǯ��+��l���	Q ��8��q$5$��+#cK�j���S�0���W���w�8���1�3��2o1�Yޛ����1ge��ѣ���J'����������e�����9�s��O����g�}�(q�o(+����&q�J��'bѺ8	2	lTٍ���g��!��*筃� t 0Ph�MH𽀲J��H(�4�#��؎�m���@��ynx�����w�>��s��Q�h�[�J�x��a�l��R��X� WV�i��J���- �5Gp;�8!;ڮ%!�՜D�9`0s�5�D�����CN�~�H��r�j&R\�7`M�-���MH��	���s��+���S�IH�8n�У��fd��Mk�i�3\�3
 ?L�F�/_&Wr*��t;�X��'��;�n��_ſl��U��>u�� B,gV+���+���>q�d� jؼ�U��f~��JO�4�tz�1L��@N�#N����V��;���@��	��
 �š���xm+ �Q��Y�����A�hv��1@�%�_�4��lO�%x�Y_>��kǹ0��!p����5���2`mH��$�d�{�L}`�ʗHm������䟽x��"����Ea���&�F�GH�z=&����n��F9�Pښ�
N�;m��e߱����*�m4(�~�j�"7m+�'�7���Y+��'))䙒s� �R�I����ѱ��Ō��&�&h��l rTj���ȸz`�e�t�ϦtBH��+�d"j��Fa��({��$���A�R��
&9F�bt�����S�w��F��1�nd.�wR�|�z�R�K�������
��^��������`ϙDK�3�Q���;pS���w��;G/�C���5Y���V؉�ϻ���g֯��n��c��-M:.�;;�b�b�����Z2�m,O�*�D��,��E?��:t~#�*�r�U0��n�+>�K��������x޽4I�_���-��1��>5��x��2a����t�2ҭp,��m���A�'l�fa1�T%'ž�Q⡠%]���n��F�/,��=(��1A�7|"E?�R�9�{���.��C�Z�bf�[�.x4!E1��Z�V9�������:Fj#��q_�/�Q��5r����js�c����aY|A�:�}bd�Wك���&�'��s�ҹت�����5���}^b�����ۈ��$�a֒�\��d)�K]s�Y�X{b[HG��+�)�8�ȟ�cdL4�W��P'A�=D�0+��A� I����Wp$�J��®�Pڃ(��b��Ы;���hg��ބY;�mXN�B6�w��4,���6�q}��Va[$$EњF��j�S�Ϙ���N��3�ilH���	&�����ɻ-�i��,�W�N��S��9Ѩ%�ξ(T80Z`^A�!A7$�C�n��j�iԑ9���1�M�Jm���$d��Dw�H/����7����,�7�8���s}~$�2�0,��<�qC��G��%�:��]���Y�.��b=����?�C�<���]�	D�`"�fh-5O6z���FB{�ࣣS�E�w��w�6ē<��Hdp�Lː��Ԇ��s��Z������)?�Q{�Y&p�M��CԝA�Sח��\��O��EClK�Б@��z�O�~�/A26+(D/"��J��F�A��JT*=.�'�m�W���v����|�Cޑ��5�պ��"�Ƙ���Ϸ�ƹ˟/�&����h^Ҟ���DMK6L��^i%#�6���},��6���w7�{�cJ�t���v�]xp�������z�Z�D�G�@UaWs��s.��q���>w5��hh�&,�tR�!��l���9$�c���F����=Jg	���\��MP�	1qt;O�I��u �(��6N���4k�U|Z����q�z����&<�Ҟ�w�����l���A��������,_\�m�u��Yb�Q�L�J�k�pI\�-�z.���D8��~w>�T��T̴�m��t�#��ֺ�@�PH�d�d�_.[��

w֡*6`�KXrP��T�um*��,;CC�5�m�%j�g���TK@�4�� �@m�����i�NJ��Q�|�޹�o������0;#r;��E&,T�P_?�9jl/�Pp�S�~Y���c�m�/jq0ǆ��V[���nt���Q�h�s�A"ne�?�:� 7�y--��=���sT��4AxuP�TZ�]� �N���A�e��bL0�`3�V^NcIį��a��L8 O 昇�.b �j|��QY=�����G����%���؏X��M'o]�]��%*U{�P�
�U뗞�'�K�9!�,�p@�0W�b�t��m}k��c}�@d�j����kK�(�˒c����*=�>G���\8 W��,��\`��"Q����u{�ˌ�FM��,V�Y�Kk�y���G�(�#�������{H��Z-2�"��_�s}�䎝2�_�˻�'p�X��
'
����@��-Ivp��P�+]������M�X�6�#aY��~�j����)�R�c��7*��\��m���	\><����ײ�B��0����SJ�>,3�%r�c�]ȣ7&ʴz������ͬ2d$��&cs<��ד�C�ͣ��I�Yu{��y�f_�G� �����"4XY.��Z����-{�Ս���Yv�����Lx��mQ��4ǉR������BI���I����U��y��8g	��c�_�>s�X2�A��̜mfŃ�U�Ƒp,z'!vNkbTg�e_M�Y��Q�x��蛛>���̒h�
]]r�"�@r+��rt�!gd�1]�� w�!����t���NK��w%@2�6������w8��u]��m�?�q��� ��G���uS��'
.�<������E*���5f�rJk�D��)�N��؆L>�J"�4H���f��^���
�4�Ro{ver >Syi���Z4��]!��y�(R�Cg����5������˔�e�/x\�Ht.�������(�@�~g�3��� O!�]
�B��p���If����q>��]"31�T��kW�8T��]�OE�k�O<�A�kB�$��]��׿��x�m�uCrG��PrC�g�N �?�}�w�����D�	ѐ��G=��z��Sr�8�T_��{�X�)n����˲���N�$��?s�:����/�c�����C����fSһ�B �ͨ��nO.��_/��W����̓I8bT�S��+S�D������Ko���ߝ�<��U1]BN���y�1��շ�+XlY��yS$�Fۥ���)g�@qSa7ɯ3i�����Rʅ@r���Ea�C"����I���8�	G./���ԭb��Q���f�:����av�z�@ܥpW��~Q�#tX���U�RʳD>|y���7���]!��-�D�k]��&�ݜ�N�{���Q+��>�	�jİ1��?����j.`	����c�پ
��u��֑~��K�S�B�e�7�薮�ۿT�2���m�6�bA�`�Q��PN/B���<�L�Rˀ�ϥ�|���R=wg��@��ES��\�$G���F�!z�р��JPF����D��č���q�J����y����-N�A����y�P/K�iE<U��#�Zް=�޺?��G~�:J���(nfG�l�EY����	����V2�Y�խ$�?ԯQ��1I� �[������~G�"�8�����T���o�植
ȉ�;՘4o\ʳ��i�fOf��N�Q���}�����0:�6�ʵ�`ngm�E��`а��WDj�K��!Ǌ!����Km\��H 2�������<�h{,��=����)���ӂS}ㅰ>I]pb�d��`B�0�g	�#�^�k\�4�Go	k�T%N����jX�߾*]G8�B�B�FD�;�÷7�<DQ:���$,T��iQ���i��(�+!�tr~�hCO�T�6����R�	�y�*�y^��-�$Y񓏻_������DEaXr��Sx�G�=z�ph���1j�p�����|�*[�u3y\�a��-�0k�u�R�\y
����Tн��[8/љ�q��/�T��}����;��� [��]e�)sST�_�g�I�������J��!n�2�s\芾��*������!r(��x����u��l�>��5�����^��˶��Lb�����l��<@�V��gP�;8F,�!:.�������p+A�2��C�0�~}�R-W�c�T6�
����I�\���C���w�'������͇�wa�ǎ���>�&�l��Ue.��!��Z�X�12y���U��?moF?��qԚ�uV/��f�j�g՞#��a0�8ֲYAb��zgQŲ#���P�1e��g1yT��&��;�*�������P��mq)�@��ʦ(8�O��6���	@�Z�7�g̋��v.�c?�� nmv�?)z_^'T��I��q������bL�%nz&+s�YR;_��эeZ�Ҏt�ӯ\�re@���l�_'�l,�hJST�wPԮ���t���'-#��;@��]��İBsĐ�����wR��_�5�8���tds]�v�2�����dh�Ɖ쬃�I����,3f
H�����p7���(sI� �Z�׻zV2i���� )w�d��Ӑd�#��7߃b��6�:�P�uMkSܼX�81�3�Uxy*Lg�R��|z.Ӥ���Ml����;&O,M�`��W)Y���R%��.V�.�b&��Y"
�v�zt^[Փs�n��Ͼ�#��=���.��
|��,�M�[������[hqs�w˵o߾�Mo�e�ƻ�P]=�j���-�P?Ll�U	��N�=����	�u�����Тh5�D����]#ue� �O����Ku�+�4oʖ[��V�E�'�Tw� /�,t��u7��5�Ơ���빎�Y,v��'e�z���n��{I�7��V<����w��)W�'-�:+�0��Be�fb3��Y[���/�����.������n���l��w]��=d�¾ AϾu�z-R�J�KҊ�oTLU�A0����J<��'�d����,��|���q�JDH;Tu���t�I���q�iӤF�
���h	Σ�o�\W[�͈ �Z�&���1F�`�r�Y���i{���y R��q�&J�)����/�7�B�K�:q�f!��K�WrE��i��!؋�� �'qyN��uH�������w$Oc���%O���LV����0X�SP(�7I��&Ë<���Q:�n8�b�fū���w����Jw2��'�td�.���iŠ��� X�P3��f���oai�� J~�v�]����?'dX�(�S9N�V�@�%��Ai�l�]z}16���
p�p���L¶ ؏����x�W<emus�Ŏ�bpN���N��R6穗����uxx`*�˖����byM6*������m��0��^<� g)�[�bT�,9_�?��wo���3�2�`�K���e�r)`��(n�R��.es�B����𨫶����}����|��*TzY�"?e�fB.oe���$��#eE1$�M��|U�ilR,�YO�a������+V���k^*��c�z�z*<r%�
�E:�[��!D{J��������zP֝�'��.�ƀ4	7��bI1�s>[n������p�wō� �H$�nF(�]@�rx���f�"�8K��Q���f Nxxe�H�d�{V5̋ �l]��&���VǂPE�Nڣ�Mg!��@2�x *0~��]�,��`x�l��y��g5�����J�� �c ;�����%�7l��M�i=�1
/���Ҩ�Ś�o��K�����AIT�pf�P��|Jz慸�j�𩧹?+=|Ӑ�@��:t"W��Z�f[���_�^���#�Z��g���P�^�=��*��l�a�]0�O����J�kg1 u!�k��#����-u�tp���D��V�J�����,n�����L B+Vj�">Q��Iy��hT+3q���ؗZ���iΌ2��h���ߣm�L|c��娈Mр�[X��!/H�!3�,mmC�RKڿ��sǾL9;���\�kT;�m��	��C���L�7!��rwA���^��U���xV���R�cu;j|O�-<G;���o�=�� �{�؄��P���t3r쉎�4��QI|�4f�A�v ZY,�.����(��P�3/0������q�p"�w��^g���D+�1��3�9uo�I8�*(�!��I���=W>�5Y*�O�ro;j�h|�����-<)ޤ�T ����K�*>p��~���y�۱\�%�i5ƙ1�V�z"'Ġ�@|0���喊�����B�^��ʷNp6�h��D�?7�f�d�T���5��%��W)�䮀Q�iub%���㪤��v�����yhɭQү²��kJ�������S[lB�O/y�(����؎G0�����8J`����ޒ8��J�)��A~��܇��� �;�$�!W��R�2f�g�02��6A���:#����B޷�Lx�fqh<��i��&1X��:;�fs����$3y�j�ә��,Bt��[���e�F�8��s!�zf;	��}d��Ų�-m��-<������`s����2k���u����D���M��%���:�h�ߒ��a&����X)�L#^X"�a��!�r��R�o:�J�L���am��z%�=\���(^K�6)�ܯnVF�ݳ%�(���%V���F�|_Pղ�^jO��������s���
v�&��.3�Ldv�9(Թy��RA����q�=L����j�H��Ö8�����T���"N���k������UMҁ���q�|��.DN�������5��Q�ϖ�X����Ne�"f'֭�}cV���+��L�� )���jl�R��E���8E�9rO4�h�fr*��4�Q�26�Q�I��o3���o��jD�$���J��j�@y��=K\+�Y�t�?;'*C�DMPd�HIgq�c����ɲs��i,�=�xw����	��t��
�Eɪ�1D{1h� H�W1J���n��7����.�������`��b�:�lM^X���"J���s}oEc���q7�7՞�U���q��+�3����r�v9�N]a��^~
��#C��J%F�!�ο7d��X�-���,�7�o�-;��<���7I�D��^}���h`����3�w�KRQ2����J�o\��W�_�ׄ�r�GxL�MI��7��%��S��(��m���9�
i�E�%w���#JI.��x6M�'̡�c+�]Q�7�p�ZQ��`u8�0��J�l��\�+e0������Q�a��5��[[?�#�^Y�C�M��
>SQX�����N��~����z�ޞ�)���8�ud/JP8�� ��mA�q�U]r^m��U��)�V�_4 �/ba�kY���H��r�Z;���o4d��jT��U�Q
;���O�-�:����fL���}�H��W����J(����B����l9�_4X�ǯ^��d7}ed��W)���YM�K�c/X� y����"��T	"�n�_E�t/F'2�z�ݦw�p��V��|$���j~"�����2U�Ay���Ny*K�g��9}����fuXf;�;��f�����9i���5)�`i�O��?�+U��9��[��P����*����2Vg���W+`d�y}߄�t�W0�B� ����\��)/�&/��0�\:��|�-�Q]�X��Û���"��M��p���9?�3�E�%Py�	����D����ҐFm��m�x�⬥��O�R9P�\�$�|MD�S�9u��R����@f�=��L���Ӭ(�`�Vܘ{[�4� za�
@�R7�_�|Y[m����,k�����h@
{���3��k���K�V�PI��F�O&*���P�)�,H��X���mt�=���L�e��j~��U�g�\����[�����ˉ����5���˒���j����tJ���g�u��q��c�ɱy��b��g��4��|�4{P12����0��{�S�����+mQ�ٯ�6�{�ٝH3s^Փy(���
�&W(���
&����r�~�Ovbr��}�� yek�أ���6>Z�h�f3"��J�!4�Y���&5>�\0�:E�4ɇ�X�&���Q�t�頎a��r����s�TH��^J�Oo�
Z��C�M�v�`U{zt�&�����>����"���T�����f��ʫ�EM��^m��^�!(�-l��p	��w�lF��@P9l�v�^H��¯��k�a�����CWz�7[���A�No>��Ko��-���v���rM��m�ڈ�֟Q,��&��OK���Ls��&���&DV���9<�p+�k�t�6�&���_���� ��Y��A�U�n���?Ԥ��,�8����=��'�7��Q������P��K��7��������[���c���n�Tb�'TP��V�Ss����(������MG�	��ȩ��8''i��9��q*�T�:_�5��������̗&Up�uU�^9~l�V[�ϼ��8��Y�_p�R�e�����sJ��-�c��-�D�?.\�����\kR �T*�!�ꗴ�����������v���Q��*'�Bc��*��\{O��[�)�c����׉\�-z���8��ؐ�y��Z󞏻G��U���:QgnH�����,��. ��_���Oq���Ի��Ӏ]"Htk�uqPE�c3f��`K�(�"Y
�G���� n���}�֮��(�c�$J�5���ڗǯ��a��8�s�KMS��W�U�=r1El_�y\1���~[GOsz���o�w�\�`_E��/�'��fv��C�F�
���L�#�$,_�$��������5m�;����m�z�|zNW�I���S`yq������',ln]�;[�P�K�3Ox��}�����'0����=q/�bJ��5�o^�	���,�D�>v��ߜj�d݈\�(~��㟵f�8AWtr��������a�W3e6M��������^A��A�5&���i�Ӏ�^�K��U`�:�Z�M�R�ڲ2Q��bb(XkI h�g�MeN�i��^H�I��\F�.�����	g[������~���sM�@kM-�dX�*�f��*����bb��@_��һ��Gh���M*)u��X�p	UYp-�=#�!PC�0�üǭ^H���1vAA��H��Jj)�eb9�W���}��C�n�sg�1�_;�<_.CKD~U�'�1���'��e���q㆐�/4��1
�hw`(;M�[���r�x�Cw�:�Ȼ�B�@vV�ۮ���pN��V�.��G��J����B3�����*��ӠE��޵����\��M����7���N���*��)��,)D���'Qއ�Ľ����A(s�S�4h���X�NcL�%�[������������9,c�V�ʘ֏-�"?v�ݝa�~�Rƚ�B)��6X�~@h�!���ѹX�������t/�)�^�ڃ�j��s��P��7��jo�3Kj��nU+��`@��b~�ٱ�/*�`��3��{ ��ZDN�Z�	%����-�9����fmx�!�x�	��j�Մ��H!�٩R����9Iv�T�)v�'���{� �6����Eb��*��]��;R`!C��~��
k���H��+��nW�b��>����󔜄�?D	��M�,#�7s�=�<��
�2��-��i�V=�ͽ=�s����+��f=QB���:�(ب�K�E�)��p��8e����G�v���*~
��I�C��~�/�q��qT!%�Y5M:g��DdԆ���^%UiK�Iɋ��x�������&�6�Ēe�����\�)��'sx��_����܇b0��>�](zb��Y�^���1�w*�qc���M�P�Eo�iP�3#�[Aa�X�����֨����b�(�a=�)M_�⟺�jA}⁾9�����b�P�^�R�����ɞ2Uo�9e&��(̜�j�����fI�n��G�GB&~3;�1"�W+�*�'�yc�$q��+�o.|)wa��D�4[���I��~�Rc#� T�Z\�x�_`;���%�8mv;����r~���WI.�ù&$J�3,	
� ����O 18x���i��չρ�H��i��m��/�۴�N���k�������[��F��{)�ѦS�;Ş8���O���ٿof�U�:�^�z��g����Q��d �M�P�	̻ ŗO`����e��+�V ���F�V��Sg0�ΩW��X�����;�7��?G.��dz�D���N#&m��O�D2$2$�r�ܵd��%�1W���
�T_{��--�|����	q5GܶT���(h�")(t7�!��$��f�H����fY���,:�����<Y�L�d�Z��� ���֡�A��4��W�t
AZ����V�<n��:����Q���R�[*�EE�D�G�'�)�`>��}�0l\�B�6x<J��(�Q]Os|��ɀ��tȔN ާ��K�uV�:Z�mt��ؓW�z���ƺ
D@��� ��,��^���?Y�즪�9V�:��'�-ک7l&i� b [��؆�*�"����}px�C��(w6:�\'>�=��|��@�u�^�{�X}�Y
Pc�Q�hޟa��77%B���n�g,�j[��.�ᗲ���u��7��`���r���[Wc���Ek7�=��g�vP�VF	3�Ɣt�������+�j^:�*����]=�Җ�Ϣ�:�� M�B��9GtI����Tp��L�o/؂�0���ƽ����{��|G9v��I����d!���'k�����pݾ�kk�c�F2 �y�ڴ���/ސ*S���=��a���y� WƲ�l�S�]�J����|�ΠHYL����?s�Y�n|kY�|���`�͎����Ѐ����$`$h��Y;i�u�	f<�*�̀Q-^� ���x���H��ىݬ�ݩPV$?�	p�)qs5 r�оo��z�_�5�z��=�a�
�_O,}8�,�
���Wׁ7C�l������������4?���Xni/�)���I�:�{5��_KA,,*�j���u�ۗܘY�T�f`P��)��� ��j����pJ����1�EbX|%���*\|�֝���3j���j�����掎
��0���xR�>��&�� n��5�lU
H��k���a'I�����J��u��!�l�}��F�teoɛ��۰֭��6��
2���C��9Q���HK��j�AϹ�?�sr?�=v�:y��7+�𔬾f�>������0�58��{ﬣ8�h��8�K�v�B��ʐ������O;��oo��A5F<ڸ���F=�:�ƴM���,{(�UA���$1+�����iɵ*�iPg�,�t]��zE��7��ș���te'd�a{+���R�	��f�+e�#!	\��|��ߙՔ?��u�v�4�F�o��7#�#k�ɗ<�Q��ѥ{ðp�����#��\��m�1���[��J&[����(���5�:���������0�'';��d��+3,yK�E���_d��Q<m�|2Xc�����ڡ�_K�ʝh����fcm+��o�l��
�"��3�bĴ�H7�L@k�Au�S~�Z3bepTrBN'�(z��>�F���G	��j|�(9�=���
�;1���C�'��1�{U���8e����1����Nk�ً'`(f6�	�2���Ԥ�k`ֶ0ZR�oȬ��Y|!�� R{����lNu�
b��J�7��+�hܿǙ�Bm�=LXR��YR�X+ŝW�nu���X]��$�7*�O�Q�&	��a��!u�ɼ�F�� R��A�� /���Mf��S����8W|���ے��W��#�/V�mK��7���~c܊,�؃k��S�j��%����U�.���~+4v ̺�|�I���N�)��gs�0p�����ȹ��F�X�//���������������!)oS���Y�I����Ɩ��y;�d�r��V�L�wK;���S�j-udZ0ڷ�R��F^�eH����I>�'��V����"���,$~�\(�l��C�Nj5)~��Z�0"����@Q��qw��buz��ђ�2t�S��-����Z���'Պ��*k�U%lQ0�9]� 4+dh7�JޝP�9{	w��iI��YO���V=V�1���?��3Dy�?"�z��%��'
�#|uut��w�¡������ ��86�U!�^��"�3��6���7��7!�?���ܟ�_�p}�k�׏�4Qۉv�+?�=
x{�;鯿��`K
p4�1���Ɛthն��VJ�f$\nv��@�"f9�6+����Tn]_8U"��- ���zv����>�C��CRL���Ţ�Hg^��z�� �xjD����Q�x�}S�#�^�x�� N�a;�s;̲�	�qf��������Y��gU@�j3|���xI�yf��\��Õ�X:�
���#�&I�+h06|y�o�`���)*'#2l�Fh���O���nMb��OTY�N�8��i�q�a$Cϫ�|���<��	���]C��M���7���xV���n3�r��V��Ԉu`��4��w˅Q��	+��-�49�]lG�8k]�<Hm�un�Q2���PpT�>�~��2���>C%��G*�X�ޯ�����>2?�X� �y��I�>�>�]<䪬cl��_�MS�⨦��ZU-5?wW�7�99�WDpV� P��C�bQ�~��%�Fط;�����<�Ų'��u��8"s�x��3v0�˵Z ��V���Q��V$�+ �~X����9�[�[���v���2
���s�<aM݌�35�S�C���ӡ�xl�0N��x5h�f�_�U�C-Pt��W�b�Bu�K�w"cU���9�B�LǷ��R۠�}Wx�լ@d��w~PK!~�,y@Ԋ�d�
X� �&j(.b��'�]"��$�%��MȱHgi����/���moو�͏�:���?��#mɽ�kH�x.��lܰ .��w���`���q,Hi�><�v��J&`�O{ʓ�h��`(�FIm�ѧ��Kj%>���~�t���RW�������%U��į+~�c�Z�%�4��-��2|�z��Ā�=[���@U��phd�����0���Y�$��bj�Y_�R��bG�3�6�9�mNĊ�𮜁GF���7� ��&C���>G6��}"��+�\� �d��>��[�Z5hH�81��ui]l��v�C΍�1��̨���9��`SI�d\�
G�h|C���õ#���û+�8�lW��v�6U ��a?���b9#��H�%�.W��#��mg��ZQ��w���r!�U�s*���V!���#�C�r��롏8�kSd�v�a��w�� �jp@h?ЂOd�;��-�;����6ICw�@]���/L�
�o�d�o�ִ��2j+�#^�iz�L	���;9.�E�J�۾Q�;5LE��B>�����pl�M������f�����X/0�t+
W[Cϯ�E�h��"b�l���M�0�%��O����b�â�1
KNZ�������o-�6�6팥e~�Yho�%�#���mP�xY��e��P��%�+ù���4�K�A��~�)5"�2B+8^�ǤC�|M3��?Ěj�}�_lra��+�-o4�<.$�*��pؔ�Zz�����0G��lΚ��%��DiO�Zɿ�ϱ#�[d�h�u^ �������Agy��e��%���V���{���[]>Oj	:ø���[��2j��9�T~v�~���d@ϫ���E��ڈ�/SJ�����G�,��Ϧʨ���n�~ d�pO���H��0�/�ת�>:������y64�M���9���,��g_�TJ���������|�A��^s��$ogL3>M�˭!��..9��7��Ẍ��N����zOO>�%�1)5��!ԓG-���檂=\Ʈ%�M��mX2p�7�TU:E���N���s�'�$��w'$w��-@@��pO�X4��E9���I�����q$��9 t�~;��b���Z��篔m��nX5�K�7���.��"G�.�I����!g��-�&mi;���r��ZD�~m�Wa��6܄+�
�:1P��+��y�uq_��&�Աz�ŊA�XR1Z�y���;��q��C�ܫ���T��־s�v�@zj�:���ѭI����r9�;&�DSU-��2> {�ǫ�]u� ^e�F[��IR �=��i+	|����n��@�b&R�U5�?��g�;���֘�5���蝳3�:dF8�V��'hV���і<�� h]��2�8m�K�3Y}���A���rb ��(E���|�Swi�it�l�֗y'�� ����J����/����%�>f>OY�4��m,e�����Zߺ����d����l7��L�3�j=c}�޵��h���x�;�D�a�Q�pCn��@(�77q��D��gu;�ؤ��O��s����PM��^Ĝ���%��i���hG-�C�����K5�|	{d��@A�Z�����y�noV�@�`��B�ip��Q�KP�"��UXA�n0+2v�����f�N{>j:�1��ڡA��%:�|��"�
�G1Ӽ�a>{v��M5[`�u&����&��� *�Ttk�G��Щ|�#�r��ۂ]+�G��#�s��%�6�P}�Dn8f�Q]=E��m����U�����59�J������<��R��k�������/yDy�"iC����^y{� �I��ǽ�����D��J9K+H��Z�:��!�KT�N	�ڳ�դZ���渦 ׭W�n��/6Q�t ����K��8*t��UB�>���x�
����G��Ul#=�pr�!=�B6re#Y��������s1)���U��ﮆ��(���P^��m��}�5+ԬG/�����ũv�~
�2�Z���*q�m (�e�+�Z6��|�f�ĕrF`���T#^��-�k�������Þ1�O��x�e�B��+�2M����Z5;��]  �"�M��&��v�Y�����>��P>�ؒ��`��|���BZy*��f]��}iy���̋QlHQ9V��&*���G�^�k���<f)��b��9k�*�ػ��0�.~G�i:�:��M����,��>
�Z�y����,��fk;���;w���L�<[%~�l5�t|>]nO�yq+����(��+���i�P��,'���</.�b��gh�����#�j�0�1\@Y���s|���9k޳��P1�f�p����bg�D| W�9��i荃l7��-�D��+��E�Ǜ{U/���������o^ɏ��-l�S����b^��>�9��$UL��&�]"��Ĉ�d�)����)uݛ�ɀP�"t.	у���`=�J�7e�wx�8���H��r���a�}'��\�ʣ-sL��5��8(�j��$9&$K��\��w�L�~� ߶�/F*hY�=� �-ˠ���NaS�Y��;�Շ���l���Ƒ��`S�S��=a����4�x�n���g�I� ��.M��[�g���d:[�P<z��0д�+�:5/��0�-y����yS�l���uB?�F���i�d}�QBĦT.-I�'�����>�s� ����������%R1�Y)G���e{Nx�=4��	>�+E�H����Ն7��p2=]f,��3h�w�V@�"M���5�Rd���h ����o�^�7w�{�$7�BnT��3]�f�]!�'��4ܭ=�0� zpɁ��O��:ta�k��7���;�o���ż���;���3Gv%��#F���"L&>BzF����:�·gm��	L��,H�&���738u������Ͷq:���o�ω/IG���|(6�(KdW�E% ��d��ǉ렟<+�$�iҳH�6P��#�j��T���&wQ��:~H��C���LM�}��[D�� s�JsUd��i�z����o�Ef�ܲR�)�5�D��s���e��z���?
����xd������mIXz�m�\��
$6Oh��Q 5����ș���.	����;J���*�㷬��mj$��2:��n%��D����m�Q���,�"#�Gоڀ:��pu�H1�;�G`�=��ϵOzC�/�]cU^��{*:�#T|@X���	�n������;�@��c����H(Ś�g�__���zr|��ߡ�c������CK0���X�h۸��T<	�!%�P<*��6�_IT\�7�9���Lq�T��`�/�s�Hi�7�'(����,��\�����a�cg���>�{��a�F#�C6Ƿ�MQ�W��G_�e�w)Q@�`��tfcUo$��w�uZ�m��yݪ�I�6�`�D&����b�.��MJ�hX��# �E �[�V3���Ml�1J�j���t	\t��4�.�J���/s~{��ui ���X�C�q��Z��x�$#撷�Jگ}���W�!��e�"!P S��Z �����ޱ,��U=V%@��� Jf:;~cOſ
���w@~�DF��Ty��RQ�K���Yd�a�/V�����L�R�?��?>_TX��@\���<>�3j��P�����{�����D1M���L�}�~HZs�޶t��e��ӿ�Pv2��۟2�c�x�>���uG���6�s̪�Ԕ�K�0+�H�j��~�/������W�,���t{�����@9NS<��ܗ��Ƃذ�q:14G�yBԄy�'�mhB!`�Y(��"�1�f�� ����K�<D���W��S���
�������:'�^�aٰzϽי�C\�A�!G��ؤF"�O�a�B0:4�^��G*�6�u��+C��W���-űj���Uɴ�KB�t=���,+��5g�!�e�t�2
~���Ae��hxR�m��������y.�?�;Q֗j�B�uc�U<f�RI�*���NH-{Q�1BSgT�T1�T��>EY���m5b0usE�x@�	`�T�։bHr+���`�$�4s\s������{p�"���j�M�N�Ț_Yϓ�7�+?�\��C����3t��O��}�,�f�2�F�5�#�\�������\?"�*�������^�� ���=�㝐�}��C�L�1��R	Q4A���o���t&������|�'��y�f���8|����2Fg�ܨ4��3_��Q��L!x���KZC=��w��Y�F #��)I���DuPU�a5���zc�-�JW����0��2�����K���',b�if��|os���%/�#&�C�zq�0��%��XsbF�|�!���t��0��5�?�ۥ����L��y���<�(���D2!�xP/>] �`�ਥt�\ �Z�-!�Rw��T���V
.��!� g#҈gp�M;�q|�j��4����)�|�ВD�6[�3��o9�jɿ?-V�z �������n�2�5��v�v�}s�x�6O��EMaf(�������4mn�}��_K9�CyJ��8MR�C_~NY8�o=�+�b���ڒ7�
��0{x*/�b�U�ɽ�R#�S�p��[�)���UcI���v����̬I
Ld�Y�^1jǺa���z��[e�0�������L�f &�����;��|����|cd]Q����·4@%yN�;'����ߌ`�7W��=��̐m�=�D��f�194_h����XM%DS�v�֤^�v5i�£����+hT2�%��9�G����jX2�(�hQ�=4�'�?�����ר�d�:.M����F�a��~}^���+�M�;�����:�V�	�+p5���{G�A��M�y���-��e�)`���vh�z�/����)��H���9�F��)٦4���ۿ*�� T��+`]�3��ӏC{��iUG�+^�?|ҥ{�R��+�5�#�m�fp$�?�Cn/"��HAo5�%�Mf;bR7���IH�������ARMm���.���W5�#�4���M0^�-ų\�l�N���P�,�c��X��t�I������O�<V���њ��l�����q"��(��b���	�0�)��}P����Y^rC?��3z@�2.�`%&^]u�e�QG�^����:�V�X|����b��^���ֈ<:L*��?8Μ���-����p>��v^r�������@���6��	0H�����dۗE1�x��(�<��-�ܰ��O���O����@��d�[���&~W��SLڌ�����b�������������}0�@��rR^�m��$����@|���oX��I��n�𥌜 �{�t�4���p�,��tV�`r}�]_깐�59���X����r'���kG�/R?�'�ѻ�>�F����Q�75��[:��<c�@)a2l݉:���;E�%b��(��܇��0ڮ-����,��Q��7�`��e������}%d,�$K ����Hb�5i&K~�U��+? �rRT�����2��zY����,2ݟN��ʑHZxW'6ߨM,>\F�-���堏b/7Յ��!
B����ee� ���sԧ�^�zNX��	�Ҭ��7
R��s������o$r(�I�nf��4�(�iGZ.�s5*>�3���z(�>#]�L�n���n�������X��"�E(E�Y!w���S��@8ڠx��@��h;~�h,��V�]�R��{'�kzb��)�4���JxV��<߂`>2D����v^�=Rs�Z3�aeb��{��=�~����s�A�y&]��zP	]g���L�b���G�6!m��I<�1U�j���2u>� �Zp8\,�T�f�C��ي�h�vb��=��b2s�}w���n�����E�z&�m5����%"�M?�i�1y�MEai17�DIt奃?AY݀{�ɨ*7���0�����L����g�X�g�|�%u#���O�M}���d��]#AZ�"�(�ɛ�_�]�?%¿Vv����.7_��6��]��5�J��G��Y*q��=�R�ڌ0��["����u��`�
LBu��tv��ˇ�p�W9�f[�[D��C�[c�TX~�~E��0;oW�_s

�P���e��G�f��S��j�Qe0
����PIS��Gw�cks=��%��ӵ��m���
L��'b#�����lb������^h��z0a��F8�C.0���a�@�L2�Ƀ��'���_kR����D�*�va���#Dcz1U����#
�_�h������YI�w�/��'@�X�Aʏ�q���-�
�\�2�x������ٲ�����>���g�]=�|����>��2u��R���ލ�c�}��WRUR�I_��TJܑ+r���&�@�\��!�X���Cr���rU�y���3B~V�
�ٵ�Ѻ��%ܡ/���]S|5D�\�W"�#�?�U��E�ᯊ�6,4��CT�$"D���O�h�w����$�m�F9.�KP���e���ʛJ;��\���)�J$^X:F'�;i�Z�K�o���D��LX[�z?�ĭ��$�xY�2��5�}�CR3t?bH���qh��|1U?�c�l��q+#=������l1����'�*ѹba �;�zs�#@��ߜ]W��ާ���5�8Gf�=?PɅ�.4J�OS~;�1�9JU���J�8�����5�BPf�����/���=�<�1{�O�����2�ӻ���k��S!u�C���~�[�E7Sb�_�U���X8�ϵ�i�v?�]hR� ��,�Ĵ3b��_�J5 �<�K�v��؁�t��:?�p��j�����W����n$m�״�>eI𴫀���B~���X�ټ��������p�LiD���t�g{�%u�o�h���er���jf���}�͠#�d�5��a�v;����2n�F����r˖2�uцj�t�`gJ�=�W�b�}�9�ju�_-��B1LA�6w�_gv�����vZ��p2����,��Iz��=!c �>��lc	���;��5CΟ�qQ�]������b���
J�H@�bۤ񄂥ap����^�,a�t����������Iej
�M��!����%��f��=V�.ٸxY���
e���k2�K����I��!.�c�ǹ��T8�v��o ��2����>�����) �C��r���-�w-HD���*b]�s'*1���B��^ڛ��9�����0������:5j�H�[:|b�)N2K��0j�5��A���ʓ��H7%���k"b-" p�C	���BC�2��=��J�H�~�j�b!�$_qxW�/���s*�F���C�J<̠�R)`ڇ��Dua�F��t�ń����W�v�G�΁�s�!��|�e������m�HQ�qE���l��1����os���za�3������D�Lk���m�.��Ćz�ou�X���҉O�B����C
�%�S ��Q�3��Q��Kc�V��s���)\��C.��� �����K�2&U
t�%T!���#�tji��B�u�K�J���9N�,�g���l����(~�`��
t 'sO�~�O)�f8J0k�vk5ft,��IK�״�,ف��G;� H:�ސ����=Cd��1�{@�_2�h��j����W�9r��i�	�O�k�L�4��}��>y�sN�#� 7�xQEe�:
��/���ę��|�m���C�2vx�WM��0�O���k`:�m$iT���ũ�Ѣ6�;ȝ16;��T\2�Jj��EoGr�m	G:]#�����7B��a���;�E޴�>"AKX+N�g�.�����Z_g ¦�)zj��e�R"W�z�t�ą�yT}��^���'qf��_1�ߩ��Z^A����Co��IYC�_rhZg��B�"/هH����E���������K�֜�n����ëD�>��]fW�Ϻט�Zɰ����v;�f{\���A�H�'�����wRTx~��]T���9��o���������.jn��ʉ�_Dp��/c���UP��1�s���Pɱ��2�D��<����rӚ�p���$���4*\oD�m�x�V�"���=Ir���'�����P��`!�n�:ʡ�fx�Q4P��ߖ&�>��0�(ศ�wl�+!�Q�I1D5����z�ю�p��-O��.-���N>'�7�����h#�b�A_o{�Y�uvM�<�];�a�z���u��]��~�� ;�١J��r�U*ky+f0�tC���bo��������|���SY�&�[�+@������%e�5W�K�/Tum�A��?���KSA�LN�,�h����Po|�̈7x�aV������z4����q�b⑖����d����!���(؀s�z�c��$l ��O��y
��{�)�Z`B���E�x����˚,����I��O+��-�7/?�+}�s���F]�e�3u�0��K��zt�� ���.�Vo!���s�zsY<z/���������9�Q��:�s��@X���[x��$���ȍu�fWܰ%�N��p��mP��,�cbd����̿T���k���l��)�,8��]A���ṽ��k��O�n�P�2�FI����Gԏ����%έN�h�B���]x_;׎�PvE0��枣5��ď��	M����D���(<D����/Sʩ�����ӸS?ʷ�x�P�߂��#�ǐ��A����.4�4�b���;)�������{C��i[��D��Ֆ䔧�W�=�&Ճ���v��iԹ|�y���x��$Ga7+�qb��Rm����x×�+����p�x����"�3��5}�ϕMc�OKVt���'�#�_d�RQ���p�SΜ%(b=/ŗ�w<2��ʌ����t����Z�!?�@��a/چbZ�*s;�Pε%wm�Ʊ�|�IݟB�y�q%D��*�@���
x���{�!�2gP��P��_z�oX���,u�sV��x}:啒�6����`<��_�X�_�ʧ�Q�.x�����ڬ�Y���C�oO<U%GQ�-���t����W�X���ak'��L��1=��P��-�����*�f��e@)�9p@�Q1��/R�m8����rI�Ԏ���MX�ZR2΁Q1BT�'pi�Ai|�������X����� �0��55%unD,�S�U��Y�4�[�p����܌�ϑGԘ[ ����g׆�Q��&�+l�`��E�_�7��"�z5:U!��u$b���n*���T�t�#>��~��Y�C�a�ڨ�yVۓ���H�6:�;׉�K�9܅���@�X��"0��:�ɷ��1�ɀe<	�^�խ��`�ޱ�"�
XK���6��S�j��xVIO[_qkqi���OѦ��(��C�Ee�Lz���G��I�v���T������:`��+�M7�P�,	�-|��>0�5��LǇ��� ����M��la�3��)0�t^�2&��d���\E\u�s�%zh�kz?m���pZڤ��V�z��(wC�27�Yd��f:r&�Zi=}�(�U�f?L���h�t&"
U>YA�]t��:-u��ǖrz�H�**_R_�3GG�%�d���������A����������{.�J��WDH�G�h�oοϛ��`B@�����
�1�d'�4 
+R�p��G�B�����ǎ�D�ķs^��4Ja����,�Z,��Z��D��t�bk������,@�)e��k�阯��o�K�t�����7�{c0E�k�@6�0���	��(`��z��;Jc��9��{jZ��Cã���?�H�,f]�Is���<�����߻hi���}6�wc��9�2��<�A���g����Z��m�)����`�rC�U;	�Xr�Ok���Z����TL�s�,u���V/��eƱ�n<�Ob�f��ի�lСvq�"���>���}jwΫbԗb�\�"��6���i�'�����8�l~��l�b�O��R�<2�߸L�5� T5D�6."EWߋ���qHF�<��� ?����Jc��R�|S�8��S`�>�A.]��%^c�4+��2�z-N�?�x7���N� �]'[��m��� q�SVW �"����;��nӋ���m��ǜpRiQ�ie+1�����d�=�J�N:D85�3�tX��~�@+�-�9��Oo܃��]�[+p�;č��O�6����X?ջ��2�b-X�*�/AP�����TI�P��ef�/�K�HW��3�*ԪЏ%�=���O>�eS�F��4�P�UD'V���,u)IaS큅R.#t��5���D�CB�{|E��p!/���;JP&A��,*��ӗ3��K�ȨM��f������K??vr��[v�����̙�Fk
ܐ�w�3���5�p��ץP�M���)�i��W0z��Tb���P��蛲6���D�&5�ֺ�ϛ���t�O��K0]�X[}�ւ엀�H���"��a�_ |e��X�z{�ج����:�2L�$�|>=`��43���49e����>Ӧ�����y�/ЮI�tH�T��AfUUR?F@v�3�B&������x�- �������L���A�a�!��м� ������ w&�{(���Z(B��:�Qgq�[���9,kO�y!5S�Sh��Bq�
����h�7��Ļf��@;(߆��0f�3�Ŧ@w&�U!���"�D��}�R�a8���3��Y�$�+粰^o�ߝ��/���SPo9�|�����x�0�V�ڒ#�
Mc�O��G�,�������6D.ʌ��.G*C�<���DK`�$!�CZ���� ]���E�&Hbĳ;n�)���l*b�����=g�!l<�K�j	�E�X.���4�RŝF"#X�N�X�]��"��Cs۹����`l(P����w�0�#PL$��I�^l���Hy���\w�~%��4���������o��E���E�~u��������|U[eX�$��2`
����)���H��������2z������?v1;j]���r�*V�h��Y��8��x�E��C�)��㮨~�Q��@]1a�+L�@�'Ʊ���2/1Z�
֤�V�X{<cS�Nξ��Q��]	�`c�^9Z�1��gǸ�L8X���ں�H�zT���(Ov��]0��	�t!Һ�1�y_�z2C������#���̓]�N�c]�[�~y蝎}��9��kT4B�`�AU�|cKjDb���Oj��R���sy��n������~���+��A�ҷ�b	��f��ob���܉��f��UB��q�l�@2�@�B�*86(Xa��د����ꕅ*a��|Q�	��ߎ>'9B�3���Cz�)���k�c�G ��f�WPS����;���a� B��L�,���\�������f��>�/ �!���J��/W5���Ɨ<��@��V$��
f=)�6��Y���=�p���)�N�@�Ҡ�$�K�K'��=�l&/M�^��r�A|�:LѸz� ��3`|�ԗR����� b�[ܜ�A�fWeGK}��EL}���kX�ۘ�� ����8F�#�f�S#0�'�F�����>����MbS�d���w���~[�Yk ]g�H�{g�jq��,��)ಆ�{I�;�Z�[ � ��A��69c�Y��H\߱S�ua���a�=r�FB�u¼ �����NÊ���ͷ]X*?(2�&�X"q���f�r�"�wiLP�vl��b� t�K�B�&!�#�M)nw�jR< �T��#[�) 5O7�I\�����U�D0�����9�K��H�tf'�����b\��}�1$��|��κ�+�/������ϊ�۵�@W���h�`�F����缋��5�|ٽ����u�z��4>�!YOf�J��@���5oں�bmN�e%�S�t#W~�I:
C�4�%H�iz�9���?=Y�����Y�3��̷;p�?���i	[�)��[nYՌ�݀�o6���QW��i��4�1YCiUŢ���gn�(̴���Wd�G�fQ*�����N@�v�2�톟t��!]�T_F^ߥ+z�K�H������"����y�!�*����Q��-�~6I�)�]v�G�-�̣�z���(^Ȉ��s�4� d�3�c�n武��*�p�������M	bCAD�)����+�
i#oBP��ͩ^��rѭS1�]��m)*�U,M�!���ȭ�X-^Uwjl�?�����:�G:B�,����2�r��CD?�hk���JI��,��1ͤa��w�ҮS��U(x�j�3ak)�ڋՕ�#:���p��ILh,Q<'#m�( ���������e��Ώ�H���fW��v����L�NN\V61�-QK�%����T5�l��N�W�/1D���I�|jO��g�|�&�<@��"�Ż,����w`�
���w��3鳔����ٝ�!�x<���WsHD	d� T]/
C�#�K��hėyE�����̂ĝ!�a��'9Z�>�j�iϜ�v+Vd��X� �2b�~� ^��~���
t(������@���##�c$�>���'��]ث�e+��{'�±C���2|�T�?�)_p'n�R��a���d� �kvc 7�W��'��sPл����]}[�-����1���(u�R��rF�_��w��|�YmRr2��Cϐ�0W��8�@#�֑
��fZ�^0�ħ�i���ܯ���[�L�X��`�?��;f��#E���b�'��b�9[S�"boI������7̸�5��A=������ڋ6۾�GH^��o��JX-`��D:|N��D�u��W ��� {~�-�b?%���;ͭ_�
#���AU��R��`�<�2�Q.���=���n��H��B���-j�:I�7�5�޻_��*6����e{���C})�OӨ�цEf�QL{���y7�ඬ�x��<�q��QzHJ�i`�O7X�0hC��w�bM'�>,ʙ��ͱ���c�/hC��C�[�q�;����8+ZnZ��BV.%��mP��I����K��^#�$K���7.�.C����R�����A��cm�#(��2D�%�,���I��r�����Tt	�G�=�<D����VI�Pc2��Ѿ����⾖��TnYdm�9|v]dq�K��a쪡M�r�,�������Jݺ Ǭ��m��6����p��I����%u��p`'>aw��B=EїPj�Rl���Iy��k����CTu��S�q�.�x��� ��.-�-�D�W
�ew����g��0�A���_lPcâ��V�� �^�X�͋$967��a1���5��������Z�1ɋAV0GӮ�'9k�r�u �z���!ڸ����y�O�>J&��E��Չ8�at2����
��DZH2����keh�%/zΛ�P2����H�%�!�"�;�&��XX�H����n�t6������1��>~1_���C�,7�5��>*�5���vݐ�����Ao��k��c*g`����):�#V`��wQ^��#�C���bax�_6�8K�v�*����&C�����B�� ���~��P]�՟y�fkN�,Nߞ{�溮1����9}t��h"Sdon,^G�ٷ�����-g�(Ǩ�*f^+�*�<�Jcьb�A��U��%`keA�����t��aO\֌��KG9���P�>́��:5bKO_�,����%Ǧ���P�l(rn�r4�@��g�t�a-��M�K�3�)�=c��g�P��l�30�0�������S��
��|@'&*fp�|F���d4�f ��� %cXhÃhR��{�,������aM(��V�`�B�n��K���T�`�ֿZ7�ե8F�RL���
0+�R���oE68'Xv~N#b�Ô�Q�핼4���E]	`[t����&�}R ���JS�f٬ UFJ�&�h�U����u�A{úEV/_p@�g�#�p�j��l�1a3:��@   O�E��^P�k�lM�N�䋝�΁n��ִ�%&Bq�\^,SL�|z�G�_C���;!���!B�)~��\mc8��m��g��8 
V��⬞�f��i��9Ե�J-�/;���]i��7g��~�g�Ls�.�4|K⛄�e5h�F-~ƕ��N�1�G�I$������>p�
��Z���~��g��K����e
�)2��@�d�s���R��1���]������>��{����H���;0ҋ����7�ĩ�׶fĚX��a�'�T�����%��
��"��L��\6nq�R�$��	<�m��?g[GAB� ��� ��+XɃZj����~�-��Z,G�ff�tĔ���D�4<�}�!��b"�̓FR�~���9�/��A�,�]R^��{p�w�u:��G�O�g&����,�դ|�E��Q,�ԏV�K����Ym�u����ˁe��{A�Cڏ%F}[�"���ƥ��A/o䤜Rt:�yqB�\�}���H�BoN�K7�8E�\�oe��+����Y�a����l
W{Aw��$�:�1ǀ��S���.�zM�)��H�<<���-d���ZC:�I�I��mx�e�]�[P�[m�fh���	�IҚ�m�Ml��DV��8{�����@w�_?Ȼ�.���	Td��`�8�� �O��
�ɪɄ����Gۛ��Τ7�N�3��6���x��52�4ie��=~���9W8j��Y�#��9R�>,/E�L�uP&�"d5,Q�t}���t���b�҃lmO.%W'�G{��V��=�f��۞�N'�p}Z�ܜ��s�1�]?׬��VPn�Yr�/�L�Y6K\Ұ6��1ui�.��3�.�pI�z� �V�b��p�?{ўo�$ kq3(�'c��a���'q�Ne1�u'�a�z�� �6;�y�� *�z�ٶ�#�d��+�<xCb�``��R��(�tLiTvv���Y�� �3�!'�Mf�y��"f�^��^�(�_�����֧6��i�����9cϛ_�]t5�N����i+�[䯊��7��r �A�=#.}���s_G�5��bf쿞���I�2��\O���	��"`�'}I�U�XG��I���^9ة>�����b�e"��e��i^�~��h {"QG��ƒv@i��艀�O}��ͧ}����Ȭ���O�M^�� K����ƱZ�Y��;@��~���ƨeP.�8-dO�*��;�,W	��?s�{�76Bef�ޒ����Bt�CvR�a떶]R�>6V��#�����Ͻh�:��f��"�dS
� ��I�!f���d�ֆ��ш��b�����rcO�N�d���h�����+pҸL&[\$��@�� ��ݎj`�Ad�j�ڙ��[�Й���fHYr4:�}z�����r��c߇2R"ӓ����Ń���!�A�䘡3%�s �)�Q`e�"��@{ r�����O��i{��9A�G-M1T�;����R��Y�xSa��++\��;xbݙ�J�j�߇O�3���3����Iw꤅�|#ޔg!�w8s���Q50������[#�}����gIήʧ��u�����Řf�b�"Bo��ѣ�MW��g�"fX눐R�3��d/߬� Amȃ�y���&'&ʠ-W�_�w#��q�b-�|�0�Xu���pY=:@�����T�V���=��
5���z�,Gk1O#�����b��eK�1 �XY}8%*���õ�"��I��"U$���O���g���Ɩ�u�>�-�&��қo�g�.�q	�fk�:�	�v���(�����Պ.��;��V0Z2?L���L{�������������@'�^��A"�t�͛��E��� ���?1���/�j�������uS+xV�HJ����S<�=�!G�]�%����cvd�Uʊ+����ԫ���O&ġFPA���!�v��ËE�s���;�, ��tg�2:*c��������d۶��S\�czM��_���붎U*��C~�Mw`\u+
�Q�d~"i�"(�CΗ�M��Q���ھ��>�����n��
 ��X��()	�'�!�����6J�2�mY�{Q�����Gr���So�D����y���� �jǳ;WT!�q]�G( f8����q���7o֑s��؉��&uX�#���"�ĳ���H�6>�w�2����5�6�y�>AG
K'��b%ב�0yd��on~��Z*3sd�e�4|�y�M�@���	st��lmV��h�NC;{ʀ�1O��Aʟ&��Y3��MS$h	-1ѥ*Nev՝�T�(��&�t�k,)�K˕�;u(�*N��Xj��,��9���H`�����_iht��-`c�x�kQc��7�Df��X P�WfIol;J����Ph
�u�Ů��i�[��V��kmT�����9;��j#.Yd'H_��>����"����bS�迥���Z��|�t�ńjɲ�w3�0��ay�x�}�@�h���/->sN4""�7J `�Oe��+�j��h�b`����V��.��W���ȼ�$W1�U��`����+��s�H���tm@�0�;�g��ZM�gʹ;�d�)/~!���]����̷B�1NCa���zeU�&��KG�x���NG�|3��Y����Y��^�b�GȮ^�+b��<xH��ɚ�@@j�~���9�e�M�a
��ަnUlh�r訯7��K�f�?�a?1��� �¬�67�[B�� W.[�*��1�ƌ�]U'G0�Q�_�M�}V;c�ŉ�?u�y#Bpmv z���&ő�p�F��+E�^�l�mg&�S�d"N[t�F��yi38I���%9<� F�i�ѷ񇊢*}P�c���=G|I`�r�Jȃ�M.��]X}��4�S������f6�Γ� ��Wb�����A�G�$u(��鉞���mSq͠���D�)��u{���j����Y�����A?��%�W�
O]���:�Ÿ��3R�F£�"��c^g=�,`1F&�F,�&��.!w�=_�:m�A%�Q&zΞ���'R���9o�E������_	.<Cl��i���69���{K��8\~8���S8�L��g��ѩ'e����Qi�݄�n:_��3�fp�$Q�c}Pb�̾��L�&��n�Gw畋4̥��4��غG�m��OxԄ���	���c-#�zd{kn�R��RL���+6pC��>�=ɧ񗛆�k������Lwk6�� �w���w����%�W�hj��u��^���d��$n\�Q�g��\�����9֖5�H�5vL�S/�}��Z�Z���.�i�V��,�YC#(;\� �e�->�T��؛�Vs���o)kg	s��p�{�;yՋ�'�C#��15B%,�$�Y2ӲT������ۖ>�BƢ��!��/Q/O�'���&k̏f�s��u�G5-�ih���N|���R]����f��8���/f�2xB*hŸ闎�]-C:̼�	�Dyn�s�ݖv&;�;���AY�[=���{�Dy�i�����
�O���AR`���1rg$�?珩�M���4���-X��6�}{�Sj?b1�^�h�K�����\����E�a3�˒�j�>@�hۍ�����[Z�gI&QeG�e����P"S�m���%ܜe���mV1���7�(�w����E�֍V%H�"�d���vS���@H�{.g1:����+Ui�g�F^�̨s�=��|��úpS��k_4Bں8ha��UQG��z�0U)l9׍�{"�L�ߤ��V�$�<��hEʧBI��l�1и�n|�Y��w�d���j�'ݗ�|�/��ZS��p~�YT�ޢ�1�R��|'�c����w���&PDr�l!��U1��x���U���b��,�<y�d�'c�\�8�^�h5��4s6FKN��h.��<� �,��������c���~�\�-R	H�w�ZT8�X)�V�f  � �R]�<�y�P����i��s�A����H��&ܡᇼY���LJ�`��P��p�c�LU���7�Py�	?�s��^"E#�FټV�+,G�g���Z�P��������8���
˓qL=��-���|�@�K΂�2L�O:��CVܐ�[��2��h��	~��h����䘷f�֛nf����p2��m��C+�W�d�=�Mp=ĖX�Y�.�Ҍ)�n�����_����E�b�M�HAI9��`�Cm��� =:��d�����E����£�G/w�q�5E{A	ǰ8n�^L�ÊbJt����o�1���������M��Gu���B0�U����nAnd���;��΂�K"� �9�Z����Q��#	�´1���鰫�F��&��46$���sa��g�A�w��s�a�ԛ�^�DJ>E�)e���"���>�O�NVYF9���b#.9��`藴�Z�X�|Sl�.$�~��o�Q���1�2E%��9�o���b�*���!N���̝
9�PV�Io�jm=�e�s�q�0�{���+ᤧ�w|����adBgQ��Ol{'���-�R�r��l}�)͊�U�T＾���߫��0�V��֕�r6��}�#�.��g�G��hڄ@׿����ӛ����I������J����@{ii��.(c'��F�@��U|�s��x}��v8��j�-6�n�ꂟjgլd�6��at`b��3�lmb�_.�z1��#l~]QC$7�#����?��H<�M�9�wJ%��~)Rs��Mګ���N��z�z8���~�	��sI�>�l)��jfh�Q^$%Z�@ޤ�u��8�˓8���h�1�O?	�����f3�(��T@�J���a>�8Gx�"k���LBN2��);ˡ����fx�D<��Jv�c�^KxH4���GьHP�y�C�A�>��H������|#��*5۝t�z��3["��2���\�z��K��?Ll�*���~�:��&ù
�+��Py��F0��aG����z�����Y#N���_�zۢ��{CZ�Fu����?�uJ���x;�� :j��-�[�&]T�[C�QH����Z�f(��u��Q�
/2���|'GULS������:-���1�X(!P��9`;P����Xe���F��@��-��ƭT��%��,PeP��l��Y26l����5_tϐ4�D��E���ZY��ݖ9���H8_�x%�ԎV�WK��t'	��v(�*(�����	��q��B�q�C�h����:��$�jf}�tB7a���	K�*��Q�S�f>(|�i;�pE��j0�q��fD�3��ځvS�4�\'7��K_�r�����߆�:��cfjsxmZ=_����u�E3��p�A��FR���cd{H�f��7��v��L�*<��hz!	E0���0p��a�ǗW�݇��P-$ ��cHǫt��A�b�����˳��x%.;eu�[�XQ�m:E�ٝ3iF����/��b��K���i��fT���b�jac�$��ȑ�XJ8����AK�0����Pg��6W���3�#�֝��9�� ��(���(��ԡ 7����'��5�bw�BR��.����Xa7iђ~�Y+E����^��!��7OWN��٣�-�f�(�`������{"�3�9���{��I	�Kb���~��T�Ԅ_�}����6/V\ݫyzWHK��N7�2��	�v��.I��ԉUX�v������%zo��z�O��Im�cL�������h��a�(̅-f��x�x�Xf?{� .��}y�W�[ܰb�LG�u�8�� 3�1fU��� _���ϑ]�x�b�a��V
ڛ�ϱa:t�Ϫ�-Oe�ݠ8�r�T���W��� *5��|�ո$KQs���7����A�����7�1�=���m3�T���S��	9�C4+��k"*������i��H��q�_����\فě�I�D��%�'�w�#�q��������3o��9NW%�f�0�h"�q~�AF���	!ݩh&���q���X=�N�@d�� �M \_�H.�I�k�����xƖiҸ�bF-��
�M�7���C�V-Q�/�-���	����h&y�W�^S��&)<�c��������[��*`G�����Ga����cp�^�}IW�����R"���f	n�nx96��WV+�����P�c�c@0�
�	\ɛ�GщP��-��(~��@���Rx����(�S*�^D�����_I\\O9��ϋ�m��Q`M��]+�'%| EgucVA��z��]Lx��Ԩ��)G�?#}$��[=7�D����pm�%2��������hduF����o�%��U�1�܃�;e�]����6�Mg��������
�`�����ͼ/2��Io�L,�<=��C�k�ؓ�6z��@�m��6���XᘚaeE�d�%�4��렋��B�`/c�%� ��JK܄��c�ZP�p��Z
Ɠ=ܥ�%��I�jz�+������i���q�u?��^�%�\#��5�m���*�Q-T������sט����iSBpb*��������^�F�06�cˊ�Q3��I*�Q��{]2�ց� 0m°֯����#1]ߺ3����ះb���/�y|S���R�>	���c�0қ}�r�^k���D�(��HĐ�Ծg?��&s*`$��ny[C\\��08�  ���zKo7ߵ�0<�D�<{��qǫ��ЩX|}��j�7�0�ٷ.��S��:����Z^2�X$@Ľ��ݷ"���j��H�Ἶ���<�ݐ
�;�ˉcw�tbe��OA��]�ƾ������W��W��z�6V����ݚ��^�ww]]��?Bv��7�1-+���}�}8�c�m�o�.�\6O#�!��5���.�wg7v��>˴Kx�O��a�SAa�MT���Řn�����6v��pD���X��@��l"�c+���e����8~�_��(͓|p�dLb;���l�gEV�[�Óm��	�^"�&�-�u�|��������D5)�S��)�$z�u���Q�ڌ��������h	o��f�"N�E�JBΈ�hP*����QG�;\�����H������wc#�X����w{&ɳ96�kD1V�	4	�@n|F�J9�b��)#��J�=s�k@��1�?���l��y�}OR-��SQf7�jV����=�b�K�>�N�G{��V��ErV��;"���V�҃��	�MJ0	�G��IMU����r����Ou@O�Ӄ�r1(=ֆ=h��#:�L��)�HX[��<�~ؚT0�
2í=�Z�:One[�a�R�{�ix*�:ַ�n@>�I� sp�\|\߰Z$�E_�.rE�1�
��;}7^Z��՞?�LG(�(�J;qEu�������>��
�w�����d�q0�b�p��\r�[�{u5}TE�l�?�ۣO�DR�cx3u�
�,���ا����9�P*����a7��f�w�J�'%U�v�ؐO�t9'����`U9����@J؞ʦ����7��4M$�����XJs�Ѭcb]��3�1�#��7x��u�Ho����\Z\��o��i"�<�@�~	X�W����0�R\����<��=�GdtY�c�>���{$#�b�i��H5�D4��Q��E�"���Y��P)N0���pK�n��r㭲Ԋ`�J��@׀-�ؾ�d������ih�>bR�����@T�k�% ^�I�i2|�1���p��� �����?��Ss{��F[�'�i:M����QO΂���c�F__� ]���H'��(�Ci.�֦=��.Jc9�[�0�x��>HR�p�!%�+�+V[��������S�L�v��@������Zk�9�?f4��U�.Jӕ��$꿹���Rj������(/4���R(^��0�S)�]�uf��Q����$���>�+K��ވ���$����p9�^;��]��%$��L�n}X �j����"���^�D���!����h� sa����ۆ��@^��?aZ�D�vAJ��E��}}���k�=�gJ�+�~7�X9�Q�_3�VS��`r}R�?=l���{y��;���/|	Zo��_�|�Va�mLUz����҉����W�~"���ta�H����2@Tc،:�}�����Ȝ|��U���w��\CFg�c\eڡwT��^�>i�K�:��j-R6��ӐQ�Pbx����`I���P�C��QsN��z0Z��x��cR��� :��,����8���'��aV�kC�uz�(�'�k�GK���-��<S �u�k�Ƌ�P$����!�����
�2�W�k�-Fw�	��u���{��b����������(��n�ŷ:��a ��2�ٯ1��`if�x�Y�7�!F>�"-��@�ݪa��po|�ks�`�3���`k"�9�A�PuI��+�.p�1��%)W57���^!��r��p7���RsA/d��٩�A%ߞ����aX�����Y��қ���P]���&�����B�ѯ��ej1@w-f�GǙZw��}G9�q�"H�u�� 8�Q@(�f�·�Ut�,�)!��7�yf�'=5`�x^�+�I/�w�H ��u�c�%�d���t�}l HR�-��KL��'�W�g�����(a�R?������V��jg�\Hвe�6(l�������������H����Ru�
:���E�5�`*���l��\Ra�0��i"�D3ȘvM��`73�B�cU��tO dQ*o���MH�v��қ[b��4.�a���0ZL,d���9��5�~J�Ϯ�$Amf\G��[�'n��hlI?�U^>�Cƪ�`�,�ۨ�bS��2{C��|,���k�B-OU��Ɩf��Q\JJ�m�`l��3	��&pKÝG�����$J�P�s���p�a�K��!B��p�RI��9p|�(�d���\R����ьX���խ��ڠ j�9�-W�xlZ}��*��F��0;��L��`��RF�3�=(|8�'{��jgU���6�m�lSNu��A�;�'&��,n��`4�% ������2:��5�y�r���3����yP�̘�m���^�!�
m���{˩xpR��Ί0l�_���ɷ�u�F��Rn�(�E�6��u5��"�.�X��ţ�>[�`[�'Ǐ�c6@��r�f�6Uc��9�Β�����$�)��cE T�����Y�#�G��a��(Z�RP%�Q�q��W��?��FX�m(�*}�`��˫ÖHU?���``%�S�3{M�}a�'u��>b������6e7�C�N���ִ;sc�n&!B���!U3�0X�vo���v���c�w���p�����A]k#�0��%]+�ě����+�F��39�� ��=�&�(�\3:��� �٦�&��
ŕ%{�.�i'qFL�TlS�S����S��:���0�N�]j�.�·�(M6k�q#Ƚ��9�ԦկS���}<��b��ܻ4����H�j�7=�����B���W�A5$ݾ)�U��麭vG��K�ux�k	��*��+T�L�==��$Z�S��
���pFժL׻��!ٛ�v�i�����,r|�#��A4'���>X$��� s|C\8�pi�$�}'&H���;�\��a�^pv�)���)���� ���8䱙�N�Pb����	u�奄R8�>�v��%��,��v�?�_��5��7�^+�dy�at�z�); ��Ű[u�5�S[m�B=<޹,�҆�Ep��%ME�ХQˆʝ���`MhU��o�[;x�`'X2�� ��XP����Șk~)�h��!����l�߶Ͳ<\?����y��U��P0����DP�ϱ�p�8�U��Ar���Uͱt�	�:}���mX�z)EIˑ$�����?��t�T��_=�q�S3$|#�q�/��h�l�f����L����E��ϻ�0Z}3x��F��~~�9о�ag.�pɭ+8�.��v��Q`����R\	\����({�\7�T�G(Ss�T�$�]�#��g�l�@�țڱ��wMOh���s��k2E���)�H�X��ˎ��s�E�*�
?���J�Ұ��P�2�mn�b'�bK�
�裟��X�	��[�W�Z%����:AmI�̨�c�f��u�[.�p϶2��`��5�#U��f�*�t����ʼ�s>���Q(7E��� H�KDetn�J���P�[���"}�@F����S�6J�lyҾ�L`�>xkF
��L�x�A����C�ď
kj]�����b��w
/$�<>a&Qع�߄z��^%���V�[V����!|�;�s�d�Uh��S�D�x�fex��)�����$p� @���%Y����/�v��-8�۲ttin��O����5V$l��=x�cy��G��@��cER�n��;ZOe�\P�fKj�򝂵}(�vka�h#(���B-���~�B�^��o|{��8i�wm0
��i1�a]O&/N��d.�/q
4�\?L����Lq�k2�v�"�����|���A:���ڧiwcw`5l뜍��쪨 L9J��Wp����s�g����r�\��ˎ����,^�7_#�Έ���s��5�����k��tr(Ϣ���Ϧ����S�x�V._�����:A��qU`N�k*b�wDR k���Wy4U��§mS��q�{'��	A3^��[sP݊`վ���ȦZ%Z�#�!��,��e��<�@�S﷙��Q�V��]��L.#�|�d��sL����9��f���U�w�x�{��j���R\�������NU��'Hɣc�_@q�zm�Y)H������[�f�;;� u:��7�p�댡��m7���
�ԩ�Ҧ�t���"@��T��3\Y��XQ������	��9�c׋�q�{�8���S#�����������`Sa{O�o��P���aC�X&v�~2]��|��]�������������n��m����-��P�R�AK�"yx�'e�ߠd�p���G��{fs`�~��
��R^��J*{}�E)hU���Z����=\��[��̞|	�\��[j��L�N��V������9���Y�L��D��O(����+o�/��d�ӈ5c���[	I��t/;$�c��]5N�����E���"�w��v�ذ¯��s�P%�А���&:��'�}ޓy�h��C�yU�Q����V
���62�%C�Ba���$���n�4�f�/a�q���Fn��v �\�.�4ݱ}��#�H�b���]����g�l�N��TK��v��p&g\�$^���^�.,nv�Yv�y�\w����)9;�2�x��p�nL���F/܉��F��,(�C�p\����aܸs��o�-&�����K�b�����d�J���^�uI�OtA�*�O�
wv?�Jt{�e�\͏U�KcI/�Y9ݷ��)�̔��R�f��B���(�:�j�'d����d�q`S��K`j��8ث< �?�$d���IzViPiF��������oK �� m�E�z?� ����o��0ɋڹ�2]d��m��lS �Ue��Tᚰ]U}uޱ��@Jsf��4�Fl���G��
�I�����
���Z� �np6��t0��ڹ��՘����������R�W�֪IgS�+M����`�1pv,������=r#�4�Z��zӵ=��:�dJ����ͥ'�ĵ�D���T�!�8h.��0�к`�P1	�C��O2;��C`,@e����]e���AoO�ب�0X�!�}�:kd5p0�g8��/y N\,�l�I�'���e}ȵ��U���U�:��y�X���6 P���7@��`3�%NV��*��� S8���.˙��1og��kz?f�5癢���a��1����K�1���Et�/9�݉�.�-ϫ+bK�\k	�k�ۙĬQ@�c��Y>��'�xL�	����ԃ�����I�ZA��t)��1Ӈ~��؂L��{WS�$���Yv���܉!���h����Q�?*8��=v�'���[�����}|�V1����U�*F�Ŗ�`�.Kg�q{���0ݵ��Yf-'��'��=\Ȍa�R"�����R�pQ�̡'oS_�Q��V�1p�!o�/�Cm&T�Y5����ID��2��(}����[C��֕�pwbz�P���.���x��5J�Q��ҙ�[Pa6A�0�ЄW6��Q�S:�����n�ӷ�����Q�w8�Ge&	T)��K�oU~t��V�����+VV�ϯ��}�c��~b���
�!��۷��Q�����v#��} �*п$��;�\���JM1�J㢢#n�s�#-<9�I�ʴ���|�g7yΊ��m���sw����N*C��.�ܨU7����u�oX4_YS���H1���z���h�)fL�^4�'�@�G�~L�i$�ϟ�X��[��f���e���Q�/�ǵz�]�o�*�U��^���'��_oN#|��ۃ�iS�)F���걽7P�C$��B�ʒ�c��}�5܊m�<�Mz{j�x�1���.4.Ǩd�b�MD���$�vZ�ɓ��$�=I��H����*�X�?V��¸n����-�@��(�M�t~��w�^Q�5��
�!��ecA�|�Q>�
���^h-�"/����*1��P�>{3�@��z�F��Ed�F��� 3��9&s�?L%�a�q����% /�A���"9yv6���1d�h�6P�V���u�ː��ww"��*��C�q/�'�LO:.�"Ώ��Đ(ׄ�6Z>�X�*ć^靮3U}o�̔�1���B�<˹K��j�b88IfvY�tD�D �,@���~�_u_��\����� �>����wKҗ���#73s#V)?`P�e�l�T�j"K2�#4��,������)�8#J-���k��d%lU4��J��L�R��k�'����܀��{��-�'��ǂa��x�;�ed!X1B���w�/���=�'-X&�m��]S쀷ٱ�Δk�Q��0Ͳ�\�	+��wuST�#��	�[���3�#f}�?���';����������?����X�7�K��g�M'M~hT1+A��aT2^��Q׃?���}<����_�w��Z,�3�hzŋ>u[?u�T�+:>�2 1�����r�܋�BEǒ�a�������4_/��5I:���X�����-*9�NM5��  Ҋ9��N+J������`8�U\o���O�2�3e�*,��M��@��QE/Ӊ�gF�w_���𿵈�"�D��t)5��j۫9�v�(���7���$�=ԥ)"�˭�G��;�������A	��V��ހS�w�o��J�M���l�(���>�e�0���*@���%t���b�ͯ��v&�G����	ԯ4)��X�_%S87�&�m���.�;�q���Ƈ��̤����7�MB���$���O�~!a�{|�{��E,�m�N�v����Lc��ᾛivJ�^p:��oǱ9�P���1�[�&�A��I��P��&5ߐH�O7�E߀Pwa=~�\�j��E�
)4��5�4���,&���Lx8�Cz�r�&�g�5Ow8��M�Wuo
`
�p����A����M}S/��uL(����)���w8A�t ������P���E�|x6~,�.����M����Å0��u�t4^Z�(����=,�L��9r	n$N޴=4�/.e\`K���N5'DY
��`O�s�X]2�g$��7WAƾ�U�J�Mޝ��Pk�����Fa��Q����Y�ƺ�g������®Á60WkJtT�ӎ��>��7?�](��w�#�M3Z�]T� ���8_����Ml2-�G;hZ���T~��Rܚ^!�Eߍ�Z]��: 9��o��nL�m���	���#��%G��Wl��5ʲ@�������=iXZ/Kޜ��ar:�o�b{̆�r���R%�r���`���sz��Y����h9�p˾v|6��K�������q�| Fս'�j�w�2%C��vՍr�g{MR�ȋ=e��2�t�(}�+��n&��YAji�W�ǚܔK�b�������ꒉ(~�	V�Ħ��%�|�d�N�h!�Db��>����8v�$�>�ftM��:�hKH��ݧS��Tv X�i`�v }6+҃o'��^QR�v�$�G7*���{	ox���C���NQ�A�oD`~�5�g[W���;Kݷ` >3�����Dt?���x�'���u\�O��aSVu2�X��=E��(H�z*?�N=���-���A!��|B[�]�_���*��1Ҥ�
�l�G�F�t����&���V�1���?���&x�ԑmXol��d���\?Z	&Q��W���o�w��M/���U,q_a�o�LԠ7��9��m��-^k����/�j���ߛ�&5cŕ�l���ަm�B�Vk��������gM?u�g���~�V�q	�PH�X�Q��H�*m�}B����xf����Ώ�n�L{�@����ih}~���<G���A<μ��p �u�+�i�y���@�k��4uIs�C�x-�x��r��Oc,y��d�+�G�5�&���&���WyU��V��/0藿Ω�wP&E�ʯ4y�+��/<+"���w�
͸���is{ET�	,t��Bs�wc5�z�k�H��m���ĝ����{�IOC���+s"��UEc�K�Mi��;�D�h���@9�B�1ԱpC b7Ov|�!ktm��6����!�yb�צ��l�U�{
��&ސ�T�c��vVe�U�������7���`�E��f�0!
��@=F��w���O�+F���ބ�hy�!��"i�,�-��K��R�������Si`Ɏ=CorY8IQh0�I����m���d�r�"-��`6X�j�unx����,O�y�<�@�9%�s'U�k��?�b���2s���!S�ρ�u�j���ŦiS�L����� o�`�ta�E��3*!w=G�T����v���>�WE�@�T�bD����$��/�������K��5ɰ]�!'-��r�K�9���\ySnTe��Ky^~���!�}g������n�g��$�����6���eS%�va���=�i%���D�N�߱�B���A�9�=�H�_�c,����K�QV�?��ba/l^�?Jy;ٲ
}~���څ��$ ����_�5�h�v1|-@�����0��'��s #Y�<��,��򹗙�y�Wv��r������Wd��0n���VGj�.��`���{�vϰ�^:�PǥE�,�S4��>��fd:��<]�)��	�O]ax�oM��&K.��TkIT�7f#��l�������)-"&�<�%�O��m|l�H|�1�sJ"� �/���m�m�S�p�SV�q��bcT���ց�{R/C>���*0�"�Cgd��WW�OF�|Ax݇K��-��pϫk���|��/�4��|`��ꄒ���!l�{
6E\(y]�sS���W������`i�Ҳ�h��DR?�m��
�U�v cҤ�#$�8|S�
��2Bȕ�~haLj�Q�ߘBd�G����l�=�!� �����lQ��vhy�梜(���=m�K����u�0q�
:�ٷ(��B㔻G�q�}��û25021i��muh%�������Ha�sY���W�B�����w|���7ᘮcS��ufj���A�`�^�E7��	����4[��o1t�ʇWF����A��5๻�T�rY9��xA��3�Aڊ[�PU�ЋQr�)���>.��H���K��=���8�j�wp�D-�;oV���H�;���ƚ9���X`�`���A�ݥ�5�$]���%D�J�L�������Ew/�ܷtK�L�0!'�p��y���~;���6�B�_���i���G�GF=t�����q��)�����]|��� ��老Q�ps���F��,x6�O�sq� ��a�P��f��������i���ގ��Cu?g�D�JY��'����_�'UG ˴B�%PR�pp!g
�J���hn��V)����k��<�E��h�.Q���-n�K�E1S1�g�Q}.T�9�Nb�01&&�/?�;f\�h��R���y | )n��Ԍ�ꖠ#h���3�R���MY���Q��[0Q %������ǃ@�����-�
P�S@ ~v#,1C�3�X�{{��%W6HF{�a�A���6�Û�as;����`G��e�eU&Lf]?	���V��#�]����)���RD5��Dʠ���ɼ\CĽ���j�$���𡴩�������"����؀�w��臿�Ν�ƻq��׺��C3g(�G��)����Z'�������g��1�2ni��2��ZU��+����	5k�$K/R�p����Y��cr'ۤ.��0�!�|�?�.(���_�͊��M���Y�T���9ZR���/�����1W�9��o���WzL]N���\��pm�_M�����6�tSa����?�Q�����?;p�Q�?xl�otا-�-�s�\;o��(�_�K��l��X�7���#^o�XԚ(ꁽ�[����ƜF�U|�ε��.��Sq������d�x�A�hc��y�*~��K�*�����>���>�������=c-2@Z�{���8�.�����v�o��u� (�Oz����2��B�R�t�-��� ���Pr�"�k��Ļ�!�Y-��Y��\u�;�<���>`r�YV+�.�w�'+��b�^��E�m��nx�A�3+�oN\u)�.��#P_LK9�i�Ԗ(|� Lt�"ѐ�-��Յ6��Cv��^~5��m8<`�[8 �����ͯJ�8Yw��au�L&�-���l,�0T{�{�"�����{�z;������������}��H�A�vW������.��y$�����C�	Nnr|�<�C^�_� �~At<��MwS�fG��P.�r�e�<�6-�K��A��G� eE$ŌV������C���P��s!�Lc�T��Zm\ðD���>6�%E3 �l������b&��R�	�x��~y�:ή�����\ixs����FA	�&���?,p�Ji�ñ��B-qGOz\U�3c>X6}>L�v��W��3�p;�m�5��ѧ����x_7��xa�� -�������9f�u��,�0�� �J�20=}7�ǭ���[u�%1ܑ�p\{g�Q�r��Xvk[H}���C�T�";��u�def�Ř���r�i�������5�,ⵢӫ�`�Qy�0�=��~�W ���M�5��䊁����ڏ�'iF3�uQL����(!��|�f�p��]:�:��&�0KO�o���8qd�����J5�lm8P`�����s�-g���]ϏJ[�3[;VW�ug������?�N���(�v��h��m��7�A];��'�
�|��/(���6��9�RGŪ��&��D�,��6f99|��CB���u64�5�*:��N����؄h�W�w�p�v�}t�B�1m葘U�|�5�9��b�ѫ)1��2ÿ��_ɔ�+��au��E�tW��e�\v�h�2Cz�h��4�{��s�W���M3_���]�'s�6u�B^���ۇWl�O�E��=���,�w�`�`pk�o~B8vng%G4ێ;�56Y�ċq�|���E[B�#@���ާn�M��n;Κ�#��h,��X�;������׃;C���[c��JĞ���<�/��W��oH�ܞ��n��8�^���-������|U0��cՁ��X�(���׻:Ώ���2ҲU�e�#o:�kP2f���3Z��?�@�=��.��`�V=Z�6�q���3�Xe��>��}Q��Ydk_؀��__�-׮���ql�7�_P��y�>a^5W��}�&���V������Q|fv��]�k_���X��P�`.>�3�\��aaU�âlG��Z G������x��c�\kmyAO��:'Ɵ���ǳ0���� �E��������@�1��bu�c��\�	��^cr�M����ʇ��â!�O�-P1�|,bY>��~��A@\5Ҥ�mA���ŷ�`��J�� �����7����٨�<Ȱ��(례��xn��{=ɶv��8�Nޓ��M_v"Z�&�U~FT@�Z[v�nAt[ ���&ﲙ�����k0ruOofY���p�S{���M�X��* L�4�%Z�\]R_��o�i�v����ƻ҂�M�x��h,�_�rMϑ��R&���ƜS$%x^�ۓV5��N��P�;�oV2%��ۺ���
����0}D�}���BS�p�+�e9�l��}2�g���@�O������w�|����(_��]����"-��E}�P���a��V6X��0�±�-�������XOC\�{��M}Tia�"���U����C캙�>�@3Y��B���tw(�R����k���ׂt���e�����(�N����;��Ot����;��,��j-��2t8��.�C _m�g�}in�
��G��iF���N�#ul��`D�e���c硎�t�%�.����G\�n-H��`�j����@΍�3�6$P��{$��������Lj��^�h��ymT���j"*]:aH\
"1�������I���&�9;
~H7�k�HTC$�����3�?},���$��<�M8mj�����L�ĕ��\�G��
E�=��'s�.Y�	7��P׶���Lĺo(fSƮ4�I�sN5���O{ KY�/v�P �U��OZ=O�n��A�I���v��8}� .�\�2/{��,{ȗ�|�L��0﹐�<8\p˞C�]��)��%��":Y	8��W�Q�Y6�B�RX���f�)���k�~Z�WI9�T��\"�|���Иx��x���Q�^��~f{Η�#X���w��P�����?����B"�s�!�:�t�D�R��b��`�k �`G\�Z-o�;��pƬ��Ǿ���-�`zꄬ�#���N��qn���+�/ 2������Y���b�ꪺ^wܞ��g�2?�I!��a��poV�Q;��Z���������x�yN�~�?T�����8�Do��c^�}��hq��=G&���zy��ۡ���dF+�p�Q�!&��uz�_i��;�_&�e�%��ߧ�݊B'��%���t_MH+ex���ڞk9��J��տpt�Z줗Lc���bl ?�y߈zRF�����W��M���&��F�{5u�~\��<3���̗��s�5Pa�@�t����$t��Q(<���&Z�U,2����+�,�J)0˿�{�WF��^�%faYH*�=��]�����]'ۜ�a^�k���J�:�5��G��-O���ߜ��6�&*�KDZ���(+N����0�B�$W���M(�,����f��8g��ƚ��b��w`��(;s��G�8��{�����D����6������**��Wb39F��θ����u�K"�2��|���OP`��[Ϣ�L|t�J��Sz}oLz$zAD˷{�ѽ%��Է���I�¬�q=���5~�WF{��^[}k�)@��P���H_�-����<�VYHKA�>�޺z���s�<B��G&	����+���jd�O,�S_���.7���-�d9�A���-5�a�.o�|��&���@9�񸈖(���+�M8��Ʉ褉�wrT�[C��mG��#��6ec��،�ݲ��kP�"/n���tS<�'��Kߦ9Ǳ���M�cU}��>�g��/3{̖�a����m���A��G�nZ���1D�C���I�'PKAa<lɕ=��?�,�kޕ��f\	2b�D$H3	NŦք�io3;p�#�Q��^HM�T9}JշK��݁Q������2�<N��I���Y7���E6�W�b��N�19�{���,X*�ݎ]����L2�;!�f�	N.N ���5e+p���6�G��#���(;�:3�βܛ�Ƒ�6f�n:�[Ġ`k��ۙ�?�����9<�X���%Z��i�>���G�����5���_�����v�e$�(��{��O��:��T ���ͷɊv���zK�!��1���WiEƝ�dmH�6�Øoe�M�H6�Miz՛팶��/�ISOp��|��Z�f<��U����W"��F����ɦ�q�?�����k��� 7m;�x�-�.���n�p�8��|C�bX(o7��b�0�U�&�c��A8=7��*�ga��� >��R�P��>{��lX�XA��k�%��QhVdY���`�j�
K�����?,�	ڭ$����6��'s�J`�P�QW�js�?+�%E��S�r��%��	����$6ⷅ�J���}^�����ą�#u�XTލ��a$��~��Ap<��]6V���� a_��,h�����y(�����W�&�rm�#������n��b�������������P��*+TY�c����NN+F��Z��ˈȮ���\�"]�W��G,n�(���![��*+I���dsx��M�R(�V uG�NK:����AW�>U��x�1i�L�{bλӹ�[�D����VV����I��8�,E@�#��5�G��/hH/n3��1�x#q/�3%����\��cY�g,�[�tM*��T>m���k��ـ��J�^ ?��܈GQ��pa����P��y+�<4�W��e8���1&VƤ3vX7/'qa��oQ9���5�c�(���T���S�	2�5ίa��=�܆:,{�����G����
 0�^t�\0�rv�@Lx�0�b���D$|��6���;����F�� �P�q�s)��Ƥ*˺R��z����� E"�V��q�����G�xt`+��ҧl��|�Mc��K`�E�I�R�RL�V��QQ���0b�n�`�\�`C_�/M��p+`�+l����B�=72�2 �2s旀Fu�a������<৕����vǳ���� �KBY|6�]���odwU�M�*�����+�_I�k���F��1)��p|YR�>��#$��!�8d����u���@��z����q3!��)�y��5�-mk�}6���s�U�R�������x��1�~l�8����݈�T�N��
��r�$�8ۋH�D�?;-j	�f��z��L�17Zog�]�Z��hI�K�neD��A�r��O�Y��R8�Bк� O�Ь�Qʼ��<�P���BN�^�;�e[��� ���<G�.��X�<��e��d�)���*
���0��V$�$@�!Mr/7W+��A�S�ۢ���ZOhд�	��	�M6�<��I~\0��GR���7�%��!�7��0<�$��+x��Fz#e�<R�'�<n�mT��u�)���ə��p�W��w������{���ڰ�\ol�����7�\�N�u���sr���������+g�g����㬾Aw��Ⱦ�Sk��3��m�e��o�w��f5x����A�����#RG�pڰ	�e!�����r��eb�PT��x��OS�����*����p�����JF��L��X� �X��������g��z��ܞ��gG 7wq�0�����fj�-n+Q�H%�������g{��Ҿ�X��|UT�]$`Ŝ�KQ?�M�"چ�1����4�r�Ju0�����F�^�G?��;H\���_c�%���Ű2���l�A
]�a�0r�F��^{/d����:i���a8~ײDd+;@52VA���U1_�Q�J
%|�@>��I�eS��V:uBQz�XV4ʧ�Z�s1+�iT�Y�n�v�QD��W��y�+��OHݾ�"��kҺ�D�DÇf���`�����9N%������!�U|���ޘ���%���r+`�5y+g�+�ԧ��[iE�k�:W� c���.���6>/Q�[J
b%O�}Z)N�ۍ��"rƂ���ĩ��Q�s�����T\ 6E�N�0�Q���7��,B�,�b����	*_L�J���y�b������?�7p�s�ėk�h�HyvF��K`iEA(l���mL0���T�>gî��	Gŝ ��]��$��Mà"���A���y�z-����'̃�Q�#A]B'k'��~��,)#�U�OR9��3o����Ru�b*"Pqti�i�(�4����_Pe���p8���h����ᠯN��v+6���Rl&�;W!J���V�҉E4r8��>�ep�!����
z0�0��#�p�������z�C�vF��q�@jր��n��v��F���|����8�m����
o㋒?L��￀WR��r�0v�����4��V�1h��5�r�G�@\��ܞֈ�qU.'�Q�I�
���>�,0�NF���G�kr�&}~�&|YO�K�et�b��4@�Ez#�\!������v�"d��P��Te�U:��<�����tAH��'���%�{�c�' �{T�dL�#��:!St*�`{�Lm�Jl]�!�B���׬a��K�����M��jV���~k$���j���&��wJ.�S�tfA���Q	@(\S�jC��w��3M5[�tPgr�<��_7F�
��P�lV4y�ߋ�-y,��$�?f�����Q�N�v��b�d!.r�!�V9.o$a�;��h��3�b"�Z�عR�J�1_��1潇3�q�_���
���H���B��F�GN���T�M<V$9�V.]`%�|�T2�N�|��@}*Dk���0�����x�D�^��(��3q�ٜ1:!'�p�����͎�R8�Oc����ґ���C#R���U�@ ���a�~���5Hlf��"?˱s�ѮQ�y��Y4��uRɶm{.��'b�]L��k�M���,}aq�3��9���}��+����P�#0�ê
q#H5�����A�^�����vA��I�=���K����~�3R�°��B�	����kab�ڗ�Dc.�amm�+�M��+�Ш����ih�ߔA��LH ƕ��)[ݥ7R�����R?.���P�z���u� �+eS���-���W~��D�9�R�����Ļ���"D���X�m�s��7b�Ez��ۥٟ�_A����u)�&M U�))Y�E>GM`@�����C|F�n��ֹh�(��r+�mZߨ7M�*xǭbf��!����62�^�1	Z���7O*�)2���-����P}���4|���F�L��.�C��k�.��6-CϋO+�VvʬA�Q����b�a0,y�"ҢU���N�Im�-a#���B;1sR���[���2�Pb�j�h��������� 7S���m��n������U��Y��^�}O�����&�%L�+��Q(r� �6"?yz{�<��T�u)���M�b����~����n#%"�k]��,K��Hc7�7�u�p����l^J��cx0_��9��٫�G=F��̚�����k���6�(�o�v��A�]�J�u�k��� ��L��k�����-��4�oS���w���C	�H��6h�9b����ͤ#��ۇio,�^X�����8[�K��;�	��d7����Ϫ�#�"�WXK�< �����#�J���Z�J�I�ՠU(R����1��o�3k���eZ�g&�<�����Ӻ�DA��ony��"G�����dL�Rh�BIK<[�����6<թ/���7���&��v`��0 MR��[����o͹B��u�Z<��P��a��4j�5J'����3֘������3!1b����b�Mr�W7�}.H��a?r�]����v��.m���oo`t��:]hu�dQm�R�j�?�D0�ܹ�&��+��ɘ��-"������	��@:�vZ��Wٔ����nHBhpH�P�R�g�����D�\Ge{aiQ���{���[���p��
���=��ϒ*�i�'ٳ?��8���3���@��}2*��$_��?w�ˑ�#oNB:Ԅ/���B����i�s6������#�z:��c'�F���C#Rl���[��K��$t���K3�5�^'2����B�7�sc���G�()0��p?'�!Z31w�*��e���A���L�@a�:ҸP�K6r�nMJ��0����#:`��7�]9���"n�`�����Ȋs4gR:��v2bkF;w��"9�(�"m���j�-n4ҟc�<��q��|��ք9��R9А[���b �_�Ц�{R5Ҝ�B@$e䗬w@����?��)�[*���?3k�p��m�x�>��`�Ӈ?y���|��V���
�U��/(�h����nJ�_ȅM7���<�u�'& W������K�]Iɹ ��>�d��]@0Ma���#=���ֽ��n3+� ��"����I�+�{ڻ�Odm٣���_Y 1@�_Z��ϔ���@69�K�NF��뒈x�״x�ގK�a��z9LZ�J麘�Csp��,������9��B��!������?�#0�V('^��kv����◳��<�K�sR�E8	ݧze[��){)�i�:�CA��c��p��h�fg���	�?���YmɌ���`_�T D�� ���!���P������	�OJ�c���+8�x�ߓ��Z��p��N�M	ܯ.U%���,�m��s��1�M���j����S=4w��8������Y�J/���+�N�����͢׌��cb�6$�-&����h������ᘝ�>:%/�g��fw} -�Qhڎ����k\�	0�[:�ߢ�УT�Y[-�<H�aa�a��I:�άg�(Ӗi������s5�{`�T����s�e��C�*���+/���m�B�Q.�?f0��cE%�$zau=|AQ��_Ȭ�h�w���E슳�"T�͒�,��ŕ��S�]aX(v��)(�=�ϣ��M�w�{{K�-Hò�o~"���s5s�-0�:�[�u�E:%b8i[������R�H��';t���q<����P�s&�"��Dg������޳b�U@�_�YȎl��m��(��̵ %ɽb��3��1��^��Q|z���K"E��Q��ޱ/���7`����J�3ڑ�xx�|տ�3F6�O��#�I�=̺����6s��]��(�&�b��xe��H.�+��:3 �; �ߟ3��[�fty�����P�Ьu	R��Pù-��j
IR-S��\A��K�!X�h��Dr��A�s�����W�JT���[��4uQ������Z�s�m��u����uo�5г2v3�V(��Qc7��?��*A��2t��h�<���4Y��./�Z����%������#�)�����w�UI�ǖ J0��06|�����C��s����?)ҝ>pЩ��;n��J�y
��ڱ��"�{S�vrF�2���J��\F�@w�j&����(qJ����4ۘ�Fʬ������(7�p{����W�YTt�K��͛��u�J�$�+�b�6Dt]�8h�������|����#X���c(�,��`���������bU�/��)u���@$�{������IN�Y؍V"&���Sֽ��il	\�Y�h�XղoȰ�Dmf\��Y�(/	�PXI9
:[�6{��V�kd��8��1#}�ߜUHS��[M-��<�$sa@;Dq
�tX)K��ȵJE�0E�V��>�)w�x���5dR'�hTi�4B�3�H���ސ�7�H��t|Ul֐�`j��Q�'�x��x�\�����E;u�nm�\�иD�,�5��w ��&Fe9ˮ=�I����l_�K�
3��ǩM�4X$d�t2�[��n��#qu�;��/N�๗j�;���d{X�ݓ� ����/�� �O/���+��Z��ly�}Oq�d��V5*[��'(���q]ꀆ�Dy�zM���Tȵɷ�[�6��x�� �f.�Y�L{o�%w亨��s`��4"'Po��V�
З`����s���3�����Ӻ�O5ӭ_���)1�Y�z�Q��y�>C}�V���Sy��de����*MK5�z��K��3z�ʻ���X�
���sG�@fq$<^��I�Y��P݃���XyjYn�E��ήz[�_o�̥�tD� �{O�W?����AS��uۤ*t�Qmn�ߏsz���Ģ����Ɨ쳒V�-"�"Y��8KG��h8��޺^ù-P��!��/�)�0*�Xya��h,������ �%��_k�j��_b&w�'4♗_�Tz��Y'x����+==�!~>�ס��&��Z[%T����`�o�
<�>+{�����wtY�����N��/P�gt��
�4럭� ��M�%n���'+�o���K�_����m/�AGǯb5.4���KK�aȺO��Z$����]*�qU�m�G�Q�<�'h� �K�QO�@��#h���J�����t�-CY�����R�8lՂFM��T ������7��:���DM�^b{<=�������G��Y�Tȕ��ۆV7A����mG���u? ��ʗ�$罩-g�]Uv���0�~�B��MV�x��#�C� ANQ�����l�<ͭw 8��W�R��8����L���^吾�p�T��vk�h���7	�`�����)����y���v�����"��M������[_,��br�Zm��=�p[M'	f � ؒ�x�hA��5K�DK���A����t�?0 ��)TC�l��nxZсqB\3�X�`�!KhL�lL��=��`P���	]�s˵������N{�Ո��X'^�h�-��YZ�Y��/�����T&ጾ�K.�=kI�mH��Hd5�T�eo:|��i�oh��%��>H������
���l(ވ�`wݲ������
)�I�)p�����P\O�5����xw��] ��;���M�!a�I�JZY�c�=!>� �_�g�H��g���ͱҜ3�aA0�Y<�?�IA'��l��e��-�_���n�İ�%�\/�EJ(��#;���<Q&��	
�1�E�9e�i�����;�`���<Y��l���(�U'�3x3C�G������PO����
_���nW�oFɦ�k.����k��ܯm*��D!:�p�N
}u�2w�g&�^x�_��G��s�S��N����������f��g;g�6nD�n����{��A23�^t�X�l�{�#���(�5\*'ܥe9���2���`�vp�]=��S�a]��VB�ux�;ڦ���6�HǶq�;&�+~T��`wKo,�2�#�)R��,"�����+����k�uJLb�Z4��Zo�(�$U�Q\#�n��n/��_k�6t���~�;�����FQ�����C[�;=��ս�g��j
uvIo		�e g*y���Ϋ���Ѥ�EnϮr0�FSd�=C�с��OQ�|o�|5��}��2�:�ړ�l<��M�ׅi#�
�r�{�uS�5�W�4�38u�%`3�X���m� +�+�Bsԅ<�=��\�M��T-����蜛�CI��OS85� ��e&����i��Pǡ /F����3FY��4����8`����5�x��vs*���X���2x9%+�5�,k[�S��Q����ʆCc:�Ub�:�����%�WoE�.W*-�4�W7if?.�~B	���G
��}ݚ�n�?�~,�0j�^�	�K;\Lk8���
�-��+h1j����?�����-0�b��\*���(��?j�Z�`@�FS}�W��QH��J!�2o	�'�o�I��Ȳ�)��F���%�B�z��:h	��V�t;�WG�1��F�x����,��׉{����ld^��DhP�X���=�J��h���|;�l&�旂Zvj�S��,���4���A��j�Dκ�f�� ^������JDpt�;���74���y}�{8����n	��y��f��<ؕ���[v�}_��ѐ��T?B���"z����(Xa�r�[t�??��J�Y�:�� ^�OL��\@z$�<��s���tm9���vm}�<(r�I���Ym�V��I��&^����'*��S����R� ֈ|:![�k�ǯ�J&c'v�Ѵ�xqa�M�B�~����T�yN��|��H����7����"���\�g���c�F��̿61}λ��ig�D�����́��WI+M�Ŷ~(��}�b�~�6�E<*�Ol�Ն���yÿ1�'��c����L��b�x<x����O�8��3����� ��^R�?�yv�Xr/�5����{bǒ�D�΢�e��9��L�`R�7�>4Z5V�f�?: �#�Nf��mEty׊{�����2M_h����\��@��30����m��TH�Ҧ�"Jf�mhI��΂�&V��u��O�ݐ��⌾+�J�&D�
�U8�O<�N��bω^_�m'DR҅���{�O����)��P5��5�-Fc��b�@��U��z�:��&DS2>�u�\��)*�vI�\�՗�=���S��0�O��d̥���%�vK������Y���w�pOõ��%D�(��[r����)�F�ٍg㲀�!i�S(M��]̑����O':��9����lu��t�Y��V����e��:�ũ,0Z����T ���N�����鴏Z~�]EIK.�!� VWۓ����9(� tG�}��2��V��h�{�#�(q��u��v������D�iŪ �Q�L�Yi���,cX"��b�ܙ&����޻�~�V7���LY���M�Q��?]V俷6����;�3cm��)e�׊�i:u�˦�^]ã���+E6�#��ٸ�ଏ����;��5�����\�
H\�`\P�9��-ϟ�)�����U��2�	�2?�����DC������62C��A��qM%�l��&�;�+fe�o'wtg׌��҆#�X��t
*��7�d�/r��&2#3�6���ej��O�"9���%8��u������������P���8f���� ��l�À�ʇE�vyW�p����	�кz�w>G`oAYƝH��Sƚ� ��F�%$?�5툥����\���13���T}O��t���f����aֿ�Z�M���f��;�J�X��\?U�J�L�8Y?6IW�CM��z�)��<��bV@���M��g�{)�NF�n���&~DE��%��Úmp�r8dZ���j�+;n�Z�P�{PvV�"�E"���t�1;чR�O�뻐?�j�WI��������m��[�K�_b@�Ag,�@�A#���5�c����Li�H?�`#H4�k)�c�K{�j�4��}%�w�r��=��(��M
��Y�
a`4Gp��t�RzF[f:�r(8�q��G�����Uj(�J?�T��WOw��#-}3\�1��A$�
��@��3l^�������A��MB�N��p�Y���0�O��'L����B���CLo:�Ƈ��J���_0��J�1��2j�&�û�]X��;�w� ��,��no,0>�
��3Y7�ZG�.�y�N��a��<�����Ms����gC�D�zb�����,��kL>����w�3V>�
>�gyY�+N�v�L�y�1�4� Z�����cN�Pf����i���� ����$�לC�E��hr���-xX��q�k��U���a� �}�p�4NX�/vD�|�0V���E�s5�� �=B!��pD��Ru���OI�J[����63��6N�nȏ��<��#�<��K-�K���MmOV3�9��ۤx��5��߭ml���iD��8��94���Z�Ŀ��*{h�[�wUs|�C��k�� :����k�4�~�H~�J��hm���D�ae8`"0�Ϗ%A���K1��+ﭚ�yrDhmy�K���=<aD�TyW���,�L�v�9��#���	R�-�����~/�H�搟��gUX\ا�C��dߓHp+g47lQ��7>Ok��P�[Bp����# <�����d���1�b#��� ue��S#�E�R����"i(����Mߜ�^a��N=��or8^�lUKFUp�3��k�����Bm���V� �!U||i ��o\��y���^�9����G�K��� I�r��D��
^��q��I"?d" �2�Em~8`��5�
���s��k��Sh<�N>}��0��n2�@���l��9��N �?sƈ��48K��7P�D#J��y�����s)3��/)q�=jC̯��٘h�� v��p� Z�4g̓�mg��1=Z�3Z��/��ŗϏ5.��m4����ų�3��IB�����Y�Bdq��A��$Ҏ���Q/���r:�PJ�<ߚ�I��A�l�Qt%�nJ�f���לeR��|BQR$�b$l�>[�ה�{h4LMf"$��Ks�tݝ͚?�ctci���;�����=�N����lj[i�)Z� 4�O��!��ݢ���}�s�'�1��2�����b�m��g��9�Mݍ�$�������n����0���w$����u�,�c���is@�PW���M����Y��&��Am���ޅPDA���2�ޝ1i�4:}�2|��D܌���	U�R�;�:����?��ь-�2
=͂<}l*��ၱ��欳�Z@��'�ZE\|���b&y�K
�@��A���k�b�����{"�O0tP�!���]W���:C�*�U��v�'vP��a�<�C�ʗ�C�
	��Έ �!���me�(efJ��ѐ�[Gǀ{կŅ�Hj_��l{�b�e~��.����ȿ_�B�l�fp���xA���f�����`4qg��C��B��$���z��/yE���eD�&!��}Ŕ`4Ҩ�G�Eq�\�1��%N��Q��}T��+s���q-�ި'c��9 �6
8G�
���x��G�tH��z��$�W����}��C�R.��!��PG��u�e*	%8���f(���I��3�0g�R���ʖ�v��ۻ:M
A��p]�QG���/E�iHñ��l~��	,^��|ْб'o�!���ڷi;����X���z�H+_p�t9�E�Q4�'�u<"�v�s�D
�0")��%�7['UP���c8���(�"�$O�\a`Ȳ1޴�L?�Z_it���ӳ���vH��1<��R;�#�c%ė�/{6{��ζIj�	�:{��q�|�*%�Oݔ�!�u����� <����c'�K|̾EzD扌��h����L���a�ǯ�;kQ�P<Utj�0 �^�.���\�d�;�+�t�2&��	˓�sDF����<��'��Dׄ�	8��S��B�����f`�|B����"7��8Dic�w�//w��8`H�ɩ4צ���O䉣����+��x�\f
��I�A�|�3��F��[��(�2ړx$�0�i3�"�[:�b�!����T�g�n���~����[����~��zh�i`�&<��[|f�E�J_V�4KW�x���'7�4I�L֯g``# �2[���8��w��������9@e~-���o��Ֆ���#����z�L}�m[�Zv���j�}��Q�L�	�%S�G�X�������%�(�&���@��Ź�ȁdh�X�T
���I�y�9��^��� 23�I���V]�#�w��}��S�<u�:���9�-@1���!T��H�]Q]�)Bq$P��\f@���# "7�I���F��T�����G��2ۊ�*��Z?�*��=��FA����h�����#�B��}>D�}��h�b[�ߋ]TZk�*^�^=g�7��G~OR]|�[v����q5;uy_#x��$5�X��K�������]��z�3�s���//��|HF����eK��^4��Ƴ���e���)ۚW5O�p##,�T9`�B���(M�1�ͨ�>E%�2Jmb*f�z�rg
\^��r=G�Y�ϒcK-��Ā���OwCU����r�T"A|3b��� �Q.Gf�4��nF�Cp��<����j��lP��=\
(_S��rtG�V����S{��@<���|(���N��Ra6��P����I^:���vvɔ_���҆B�!�o��DȭѸhk���y/�hy�9��(���  �W�9$�4�ރM�Ŀ/�6m�n�s�Y���E��aW:�"�Z?P۷�dr阳bZD��@��H:i���K�,]a.����,���u��/�{RU����㣦�����{����7�{]�Q�>��	`{�T y�2�S������7��~�E�)�k����pjR����*ɞpҮݣ���$M� 1B���r�x���c�zDv�8�R��G%���[dd�I��IK/�ۗL]�6�ޠ�%�Uq���!%7<�ZԢP"��H�l�1ٻ�	���r$(�KW��:nMkI�*��[W�<��!I�I1�N��R��7d�|M_Pr_��B��"��GęQ�,�Ę�JEɤ(9#{UIѭ2pH����?�u��d��!e�s^��QԱ���9˰԰r���K(�uG�&9r:U��������w�ܛ^K�ɣ��V�쾀"�R�w��7�,-*��'1SE˧a� 3c+�;�/��MV@��A���9�E���D��g�����5�I����D�=������;�P��szH�����ׄ�_��\f��zv!j�N܈FN;{$�{6em�ʼ�)����<L[Z�<gr�gbCG���_�L��f\dpO�Xd�e*�F�S�[+�$�|(ď�_2>$��%{o��T���B�4�H�䓞*Uҟ�*��<a-�gb�
)S�-}���X<�&R2fT��05�.��I`�_�@�7�oZ.���9hJ�Gy޲�BR9>?�T��(��xg��yN��9������x0Aw��4r!m��ɥ,U
�v�n�`�?q�1bR��i8��b���þ�����{X��P�:DH��<2���K��9������+��]�Fj��Uh�{άp[_����ǈ"���?�ב�\����l8(��^�u�ֿ�u'���V�٬2fz��4D�]�uYA'}l��Pf{��|{��^��`�W�0����`���e�c�đ.�/���T���
�@Y4W_��Dܦ���e�5Ҹ�"fmù��a���\����V$�N)�
a��vI7п]����7c�
����q�Lb�N[y繖���򍯾f�U�+�� �ƥ>OL������"
��A�)�*C� �R���n������x�%��m�WF��١����0�Rj}v�fɃ3��*��k�v4�F�-7��o�����<&�������p?��U�a���v/�+�_��򁾅�s�Y�G�'��o˓�Z�>U��4qKhմ�YeUl�������/�#��P��9o(�k��ed獴��O��#P�W�JUq0T��$W7��˨�ϣ~v�K�x_rV����H��!,��q�1u҃"�ٳ�|�-����îv�^K���'"�>
-D:���q�9��<R�����i$�n�8>c�.�W*����$솥���(��-����W�M�׼
��W1.%u�6}nt�m�g��#�'�;�����}{�3df��tҨ���6�r���E'��**+��F*;�t��m/�����
�v�5�ي5�}�`�}"� W��Q�:�3T0�x{���	����ZsG{T';H�#�:fߎ��.���%�9h~��c?f���ˆ�"��c� �=�@cWv�X7YԔۓ�l���y�Mr�zeq_Q�>bs �[��-��S��JH1x�_�d����J���9:M����z���'�>����mj?�eR��1�@
�E����~�QV���|�>�����^x��!�����,y\9�;_��z ЛA5�d�?�4ڏ6���ҝUi�f����$w�FEAE�Q�^���P%E�p"�*��]� �?�������5�.�+H��'���APZS��ɖH����c�su�(� �U'��/���"�G�#��H{��FK͘w*&�B�V��UǑ!����:a�?ͱ��h��г��r{�O�.�����߹¹*0�{�h>0^H��0��B�7��}���M2��.v��@�-����e�Wa��f����\�.�H��j���!�d�C��d��1ͯ��vc��d�k;���"���*|Z���K��-o��O@ϛ�D;ĻZ�^��L�z���I79\�Y5W{�j&�|�'}��S�^�� �,�b��iL�{�Ŗh�3�3A�p��'8&�l@X���YIR0s�CC�#րmM��|�ڪ=����Z�Ra��NTƢ��[]J}��x��鸫�&E�H�wĶ��l�p5-ޱE���H+R�h����	�2�ם�j2[���:V�Gi�,��e�����d]�U�m�`Ȓ[�7�oƀA62�<���QElu���,g'k{�=$p�܀v��] ���r:U������J��|v1���������7��ruʲy��W��9oVv}7��Ѳ���U55���μV/����JƓ�Zn���8s�̩��j<z� ��(;��p��[ii�6�ĵj�6
�gS��d���G��N�㧪n�?�(�6����K��D�DҢ���'g�J)�>� w\�����F��,��0=��g*avf<_ 1���G��;4Ӷ¯6#i�������kI?�.Ve�x���ǽ����2�=����?뮬��0��πs�E�U�m���7�^���8��s;N��y�!�����75^u&�'-���Mn0��;�.b/U�g��_��gm)T�N+�wh�	@X��>Yn=�i|���铼�^��� ج��p2�f@�@0�Z���eLq\��'�3�������C���mE�Q�sH������5�`����(�s=�Y���E�=���p�W6����!�iH8�K�3)/g���>F P7fܪ�p��+hi��P�N��ʏ�;��C/��m�q�jL��2��6V祾 hlռԮuq��׹(UbQ6lw5�[=�w{ln��|�jt�?l�V�+��Ňi�ۊ�yw��3M��� �.W�+�u'�Z{�"��
xs��[D�!�9�I^���qG����������Z���ɟ�o��5W���Ƨ�"���4���8�J�M�G��fr�W�z���x,5oy�1%�Y
/������B����R��yeӧ='�倿�4��ie�M��5��uce�����q�T=ɲ!���w��c U'�<D��Wwb ك�g!�Pަ.�m�)��)GKvݸ *��(�^��}�S`6�ɅE�V�e�y��6��lRG�f�B{D��c�$����=�Q���믃]� D7�%;l�fԡ�#jjϡ/1���H��k�ogÁcxK���ge3?��no�˸s����N9��<sl+�[���|p��q�5M�|!!��f�f��,S\��E9v�I�J�u��g��>4��v�0"R�e5�.o F�%t ����.p�Q�V/�j��D���ހ9Ӽn<�����/,����]S�P�J#[>��'���d��C=���h��
r$�͐�����QB>Uv�M��� �!�I�����	�o7?�L+�9䰶2WQ���8+��k�?�CE�e��i��-x=��m�!pĊ�+���Or��M�Q)eg�4=֡T�DJ�X��2~�@ӎЀ����'D��B�)g��)�]��v���{-�?g��H��0�!�;/0]��A*.+�S���><��#�uN�1�+�6C�w�A;�7���8T�"��f���^�&�Qv���͔�w|�_	�p*�����'�0q�Yj[�g򴬈W)�1t�t@G�L��6��x({�8�FOjVN��-g���%q������'�]��mi�s�?f���vz�a���ڼ��*ŉΰ+�:�|�o��2\���j�}��k`��G=bw_G#��R�n���!΅���w�l:8%����m� �_9�6�:	R>$�8�y��/��!���CFh�������R�t�!����}	��7��*�����Z�e��tZˬ���K�t��3 ��v�y_X��a|�1A3���,��r�V��EФD�W��duE%	 �A�X�'�S���0j:9�TҦ"�yh��U������_��-h��<��f1���8��,��-0�/ɢPO��%�#��������ފT�0`aa��IJk�g�<�%��uT��n�U ���u�C�I�#�I�rښ�o����iw4F�9<��P�<|u���+F�qؚ�!]���ȼ� ��G�l�v��pq5�ǫQe���
;S�4�����<�z���������	��p�2/~o��#�@��$|�7�!+W9�b��?���FUb�;�"�[�ϦFq�=]E,�<�V�7�ۺ���
1z���N�?��s����r0a�C3r����$����q��e����t7	S���:��@t����"���$%���P����==ް�;e!@���S�*YM?��&,K��)7̮Q�NJh���;R���7o�>6�rr>竛M*�!�>�wwZ��z��^^�C��"!4�
������Rƶ
3���#�,�	���0J5"�l(�q�c[��D$�
q���=E�ƛ���p6b�BtzWX~���ݰ��Vq��!�ږ�ݼ���C�3&G�cS�;�%�吧	���"�ts�}�q8��6��z����[�2J��:�(��1���r�wL<���jۇ6�[�k��15��?t%��JM�\B� 4��s�D��b =ݭ����>@@}r�O�LL���&��Dc��E��s���I@	n���p�����|Kl�gt�^*�c2�}x�4?z�DY���@`�u�׫q�e�C�h�̏�j�VK;V�KI��r������-RAl��a�s����0A�a&��I�!����U�Lc��j�yd0̓r�(���5�L"[�R|e]��~RĄ^���_�Δ�r��
�隔)����}�4�p̗Cr�p/�)h�\��,k7je �RE�v2���X���N����M�ұ�~�@�+<Dlo�nM����tG�A�5�U�ʍ׃xg�j�����/�"Z���:盿�9Tp�v�m�;{wF�߯*��t_�v;�5��r���o��]�,��� )�"m�K�mE�<=ۘQ\�>���TҀ6I�tP�}8h��<��|^b0昽{�?;���_�z���w�-�@j��?��"�	1s5�9]�L�n�Ԛ˴f�ad0��	�f�- X�����qW��gM��bh=5�zV�q�C ���{�.�߇�ǒpa޻k�Umבk�!<>���шЌ�H�B{��B�� S��#�A�DL2GH ��
�j��ms��"/;rW�b0�d� w��)8}�\w�W�oK�3�����F�����~G��ާ ��T��Rp?��׊<D�I	�D��I�xĺ�$&��ŵb�yY�n
�����<���-d_�X��q�`��x�qW��p}�i��8�!ڌ*;�q�ɇB% ���Lՠ�`�{[+U!�2m�X���[Hd�A���V2X�l_+�lR�u䇺�Z�,������d���Q}S�������!��4��V�T�]s�
b��3E-0�����$U�,�̤�/RW��g��$*�Zע�_�͟�&�kkǦnk�n��hR������g�?�)����-��,"%T�$B�ȦW�D8��~E	�sa&�����H`6�U���'�6��9���Tw���<i�3�˝,�x�L<	��ACB�g����Ȗ��e�Z�)A�~���]��	?��=�u �Fu�b,�~X)B53ʝHM��R�����fxש�@?<�	���a�	��ޒd\�JNZ�+�Ì9M@j@�b��;�b<�� �����&Y:4B6\�a�OR��2��N:�{����6o�縬z�{G��v���l#�kN#�$��-`A�S�hFh�����{��H�;%=��+�]�� 	/*�l�ML�tP��u��%�%������Q�l�r+5� 9"K.l��G�� @�㼇)��D�����u��Kwiq�������RUL`�^V�s{�Y��"�7*�͍?y9bó�CN���b	D#��5�| �IQ���x{Vr�pQ
o��,��s���"��DiO���lÃ������9�-���j��!����Nv��X�V��D4�_^J�&M�����W(��(N�_CK[k�
��C�כiF���G:��d'�W5��_-�8����5���t���s�FuAZ�_J0���_$k�fEø�u\z(�����պݼxrf�šF@��s���pg�oR H�X�=t����ed�AE�J|�r?�!�1 ��Ũ��lu��F��7Yn��	�;q֬gu�I��r�7$PJ�Az���#�ٖ!3`i�+*U�	NN�76�1z������,p��ȳ�+�*��T�)R}�����.��v �ѵV�c�~Z�b����lݤ��]ѝ�Vu}��N����������<\�"�� �/�����
��~�1Z�z!#"f=@կ��h�)��	`������}r���������/���{�h�Ѕ{"���&��R������H��L=��}A�)��P ��WaK��9߬~��j�Q��,�������9fD�5D��Š9�3�����RzN�nv�4̉Ƃc:������Bɇ�)+mg#�}� &V���(T�P����E����|bg�
����x1�[@ ���P��:��β�0P/�^���ǒ�-�ed5�G���1��O2�@�h�U����!��O �eM<շ9�,s�hǻ����2S.G�w���C���p�d|���-��d��W���`G!��U<�p1�1J����4�o ��V���!��7������.+ ���X	����0Rٽ���L��&S����g��C�g'�l���-�k�Ww��V�0r8J�X/<����<����a�Ve�
���/������;[��1��e�{�\1i2.���eǂ�i*�]�dgnߠ�VԖ)�H��NQ
��(: ���U/�!�R�?Z�_8]��aBk� �_8-�H/����@.&����E�r�
gIOя�b�Y�%"!��	a�+Q��()�ϷM��*�$޼6�W����}��	�4�q���c�����f�:�X�O�w�"Ñ�D�տ�H�,p�=T|�yQIuqt�L[s-=�_�_�jB.�x_����i;p�aȈ�:�񘩮1��1l�63�~0CS���=�6���$���}M��*t�EУ"��5d}cq^��y��بKDGY2�dlg�� CL|��lc�������N[h�x5r�6^�]�D�,.vzC�"UA�b:n~�;L�:)�؆�����|
�	<>��[3:���۞�;�b}V\��M���������?e��IP���}���^�>�e�E�T�*�>�6��	^��S'��f�I$AšS�?$������Ӫ0�	.��7EG�o½T����{��0	�*S������=g	~r󑄏H�M�?�{�&s�h#@RG����msA֕����츀']����yS��^���/�T]|@�mɿl/\*�h�N�,V�^W�ڔBϑ5�����Vg ��"Ř�3���崛����1�K�'9��N۽s���K��	�DըD��Z"ta�N���m����T�=R��2��fؕ�����6���L%��ƕ4��y�(�Џ1qeh���M"rx��^4�W乔Y-�{��]7�������f�ğqBP��NBp��G�@=��Ǟ??B�������=��'�6�յM�a���4�#z_k��P�,�Aǻ(�&�`<kqFӌL��Y̓	D�x�-X�A K]�m���l���y/C��0q�~l��|��X#�O�	�Cc�j����B̼J�䬸�C.R7�
O`�H��ē���Z����	�9��'�kOG���H���q�Ȋ�q����'�����d�)	H��}c	x>�Mi+E rU��y̯>��uT4�j՝i�%Læ[�w��P�r8�5�.�/�@c�ha]�Dj(�H�)�ZwIc�Z� ��<Ny��A�8D�6�`�o�nA�5!&���ݏ��9�����f({����8g�PӪ�*�oBJf"�)�p�~�)�gj�~Eg�@����.��g�3G�Ű<�U.�RgSP��*��̭�A3:��K�9z�EV�RW
Ur$��t�K #�����!-X�-Z���`����x
8��s��ڥlP�j�ZԤ��z��Tܚ�����2�.?g`�>�N[�Z_��=��O��BԀA�Y ��VBs��:^��"�#�y��ٖ����cgB���EDnP�5͡R�ׂ��C�)b�@~M�}4,�#%��I1����X�b�_�W�פXn�US��G��z�Z�D�q+"pH-��-v�A�T
wJ������F�jǕ�3�]�(������8{aUs *)�Q�=&C�����|+vލ��q�`��E�B6D�Y�����O3�P�)W�ȓ���w�~���⿱�D�������1~L�"6�Q8��_.Fv/q;mRR/S<̼�v#�:�����Y=&7��`����yQ!��%nM�����<�O,[`� ё��qn��]���_� Q@C�9_ĕ;�0�Ct�̓}Oq6��4����:	�X��M��<�@yFڮvɎ�����:�W
�mq:��i{h����6cP�%16��;�3�r��ɼ��ʲ���O�<�n�՜+�uE�s^��UDx��]�q�^lU%u0/^�4���օ�a*�.t<W��$MG�TJ�����@������N��rj�b˞����,�6&��&��N�0�qV�+6���_�n���y� =��J�`�Y9`�����{�6S��?��EZ�;Q<�y`;f SQ@<��R9z�<�t�eZ��2'vڟj�\'M�À_�1_�i��]�����1�cq�7�\f��`��X?�y�{�@��PP�J�l�Vd��,��7&%���U�	����J�/���&��Me`����co!��Y�&Ɯ��U@bq/?�J���
��CY�\��B`K��(kQU��y��=�헔rz�&*�;ҥ����L�!랤�/H���3���}!�E���l�*!��'�s�$�&�K��2k@�$|P���**�4�g	 H��7Yw���:79��u�J�fb^�U�#�B���b�����`�a)R���&�!�d�/Vm����} ��B֪آ�L.��xoB����&ﾣ�F(.<oT�����P���k.ֵ�M�� qjN��V�3�Fj����DW0\ٓX��#�ER�?��V��n��>S�ᝇ��P�[~7)����L�s#�\M�D��,vg���Ά"NI{\X�Z����s�j�O@�|}O��'K��Ǆ��m�<{��������-�?BQ��^� ��`�_!����q��y$K`��q�����h���\.��K��lB.uה���Z-T�8E"!׳�ްV�3�%t{���8uډ<��ΓR��Cc}У�y���{���\utM�En���I$]?Ei.����������v@����0 ��P���òZ :p2�;><��FTWb��y*c���n�~��2�R��������Qtu�̞~�O��� b_iR��dq���.�O  $Q�D$�R���;T�����څ����k/M�O{��\#��n^C�H������jR��ܰ#�.�7w?�N��M岜��n���m�9�����N��8��g�X��yº
z>�M��ω�#J�"�;'�U*�� "��ޅ���"Grd�W-Ef"z;zj�C��֑;�%S���o8������y���ZG�؎<ǡ��U���>e�^7��~��X���v�^�A�Z�~�b2l+��Mګn�����Q��Cd��kK�
��V��]	���D��-H~���v��z�R��2�ڽ�z�)u³�T�w¹l��/��"p�D~�Y�1�(r�ܬ�c�/��F�T"�2� ��C�Y���� �"WծAj���c��ή���hPۿ��:��%��[�f�(�SqH�|��p����4�Fc��N��v�K����|���[1i�qcPQE����C�I�^2z�N;��"���I6U�j��fڠ���D	����>��*�_�Y\�5.�KN^4�h�`ڹY�:��p$����MU.���spY|3��.��a1�O�����F}�+��r7q���V;�����L����<ۂ��B�Z${:�9�z0��CPt�x�&U�(Y�&(���r�W��p6�z��9�}� �ͮ�#���oV�X7�AěC{�u��&g}����9%�s�o�)"���4��
8�Vٝ��>��N�w{�U�������:\�V�B@��>/M}`�԰)��V�gj��P���ld=��w�͛Y�^�ɿ��w=טO5?X+	��h�G៰�.�.�Բe���	�\n;	>j*$�|���<�J�G�8�"'� �/�T�sE(�g��`=�� Jt�P>h*����K,q/�"��|����:�����;��h}����w����iNi��R��d��z֋D%w|�fme�u�bU�ӴO�̲l�#M�K��o$�e[����Rꛉql�@�`�攷M�͕�i�r�� v�˾��BV�ϳY|qY��ER�P�{��d4wN�.��Q��6�%�[�RG����&p�缢��K�,�q����д�O��n���:�����E�Tys*Q'u	��1�\8F���R���A&a���{֖ �!^*7;�^9�L����V����T�-"Au'�
��\C7	+��ߞ6z���=������d��ʉG���ˍ-�u����j5��v�~��lDz0N$w�C��B᝜�l��O2��Cs9�B�jw�$��y��2�g�{��v)��{r]miIWވ��"Ԫ����Ͱ+�Ǒ��
��fr݅J�@�TF4��a���حH%��ދ��O15�{R������/C_�^7�%I���bS$���Q����`�3���>�����ҿd���#�ɔ"A�zݽ+dZ��B7Ո�N����9����U0��$8�f� .���fڠ|qZb�^c���"�X� �T�,���:$�{ Q�oP></{w�U+%0�f?�`B�n��>>�m�8P��Z��n�/rˤGP(��n�&�8�sFW�Q�g_ӓ��U���7p_ɩ���1r����j��'�I���M_���8�=�0@�Rʴ���j���.ތ��GJ	������ʕ���E��3�o׮�C<&�0�5�"��H�v�N;!�E�	ʇx)����>�_Dᱻ����FƢ�rn��������A�|}DT�1=n1�=LD�ْ�>�W�H��h�f��̮-�C4/"���%�ȐX����$�����*5�O��{�G-ͦFӢ�X@}7���߶��Ay^��69C����Q60��H�w|�3�.�B�	xg2���,�/<���]������*A��G؟"3���}G1�D_i��b��;�XV`t����ͩ+�(+�,�%��u��#�A�D���y�ovD`d�ہXxx-X�nm�s�^V_�՛t�v�cc�ǃ��?i�po�~����������b����yة��g~u�o���l+G�= �[Q��A�4�Ws1K�6�5Up���.�-�PZy(��#�0�6�@avJ�aF:��!@��k�/���5#�Z$����-<�4:�غ?�9�h;���;@pr1��sݒ��9�А��v��qѪl���S����  �Z16l�-]���f���M!�]{r�?�y���W�)��ݏ4H��X�$�W��鑇����λq+vC��i>�@�x�+]�o�c_sՓ�"�+�>uޭ�m�ľ�� 6Uj����!B�-��Om��[BQG��+ �9hK׀�DL-���*zk�lQj���s�%��� ��4/�ˈ@$�6�.��g>a�7�=<a��t>�kة�	K	���֝��9�p؛%��lT�=��Q�F�����jv{�x���hhkl��^|!�+�HQ�)[���g�]��!�"i�u����H5ߕ�~�v�?���;7���u��!7��
C�h�|&o�xS:��=T� M�33�NQ�"p��n*e:m��K�_O��h��\(�����<�c�Z������$
�J��Q&���3y��a|a�LblQ#�f���Pk��v��?O0�XIH�yr�R���MYؓ�� ���\8���Y�����HL���>��霮��������&��3]GVJ�9Ċ�{U�sn����gB����WUn t)����nq�0��������sŖ�	1��fcV����EOO�ˆ�M��Aܨ���U)������^x^�whFC׆�#V��+y/A�SY��;ٹo.myn��~�0'Y�S��V�i�68?+$��D\��ޢ��3�ǝݠ���7n��ZT$��)W�/�A4FC���+C�I!��Q��Ycp��v�I��-$������M����A��/�)s�,�J�uZ!������FKޠR���V+��q���D�*�`�{b�&8C�`��ba�vC�����kؽ�Nw�6��j��W҂�\�;H<NP�y��Z��O����ۇܸ������L��v���ζ�n��r�2OZ\��A-w~��u����"����e���si�Ý���>q��k�c1UG�s������@��������o;�\p���L���l�eF�2�+TNW|�=q�ze�K9��R�����MzePt���:߈��w^nä�G*���~iI$U�y)�%��wa� ��=C���SB2�@�`��/g���O���O��"��HPݍ�o�p�;��ZA��N�_�N����IU��3���J�g�I���F.y�,n�̡	����D�Fi����1�=�f�
�X�7�ڃh3��ߍ����0I��q����%�Λ�U~�c�Fm�"�O֫�g�: ��؟n��-��}� |��ޛ�ֳ�V�%� ��A��"�y>����?�����?�ڵ�M�k�jbD������>i+���'�󆡍o�|v��;|r�Ԛ�(>j=|��Ե����ߨ��������_���[��@�@��4!m�Gi���dO��¯Ť �_�m�p�x�럠�}�)���?�!���Dt\���w>�$�n!qMp��F��7�T^	�g��M�e�.�˅T4�|��[�X��*��(�oD;��ɇ-;������U���e����ɶ/���Xh����9�.�����Id|�d�pJš��/+g��1:�<h�by�j��_�ab �f�K`r/#��Ⱦ�����7���3��f]�$ Z��!��"m�3��ۜ�%|KkW�\��|-���OQf��wp ' ��e@���JF��^:)�&m0��!�:��.e�� ��Q��XuƦ�\�kD�l�<�;����/#9��vTnJBK�Y���~�y���'��>}{�c~�HC_N���i�Zh�˓�g ݋�̯gK%�kM깩PF���*8 ?��9f�N�Ff��N��q+��=oF�/�����`o]�Q)�cV!al�+"uS�Ӭj ����1NB	�����[�Mc4 Dk�H��%�l0>�WV�ge�a2��7vmk����]�]+�K	ǭq,0�P�F�JjU�	3�!�~�7�K��7�{~Q����@\��|L�H(k����B�v�Bѵq6�(��7P�<��@Z�	{7+dQz}�L{y6ufF��}CR/�W����2�n�qB%|�b��9~�J���G��^�v�CI,*l��PZA���1��R�Ge�QO���^���f��:r���/T�)r`2_c�FÎ�M��;#6C��%nY�K#���1Ĵ�j���s�v<�[�H��?�[���5���-4��8�u�Ih���Jk�m���)�'z��^�M��{��u��y�V��!���_�]�h<ޅ��@
���|�;�U���q�;��-?��k���DI��M��B�9Ў4K y��
�K$�ET��4em�Xh����&
����t�Jg;]U�1���q�����I���������0	�V���W$Y�C�D��u�p��a�WV#�yO-$�V@�T3�ZIX��� o!�H��7cw�$=�tc�ꫬ��I4���g!�v�H��3V�de��3;Y�x����3���� �	ԟ%��yF����k'�^J��Gˉ����B��M~v�=�q��ڏ^�-W}�d�Xm����l�=}Q��%�7Pv�,_k"�BD�� ��yd�#y�d�i���m
:z]J���A�i�b���!�Vږ8Ʋ4�$�
J,F"��/�=��{W�$�����굲�ޠ`Yg�f�%Qa�G��<����C �6��.����|�^�y��	

�������~�MV̀Ը]��";��dc/W�kk���M��K!ei���;��k/"�R��*��xk�2�+�H�O$���^��k6Lij�K�2��sq�,��#��l���K+�������)�}�ŵC�y1皖_�W���ޭ�M�3F�&I�T�W���:�i���'���?�`��݄<YWC��t�<�7mX���B�;'�ý�g
?�p���V(�4ѹ2V %�+?�ge�pv��N��&�[�B+V�4�q�����v},"1:�!3�̻%�4�����x���6ċ�s7($��R%�?�^�g�)E���_�r#�[*�i�
!���*�9Y���vs��q3��4��G��*��ܤ��G�޿�T���3{����V�	s�V�ư�7�S�q 	9�x�>B~3��Y�6��.�p��ϒ|E0�ޯ��S�飫��0�ic/do���W����t���hm%Z�<��#\90NQ�=�ؼ�^,}C̽��o�?vhg�!n�|an*$j��,���Ȩ�b{t�S^B�h�yA ��M?f�7}V���y�1�߫�/fe�\��g�S�l�<E��6�v��o���|����!���{C���z	5���Ot��5��,�EK�D�1��I'$&M+Sv�l���8x�ʱ�d-�PH��D�ӘY�>_�y.,�!v���X�z���P7�x��$<0�����:t�
����*wr�I:}�db8(z���1�S��+��ѐ�Ԩ`V�1�8�!�1'#��!7�$o����U�Y7�Tv��ϱ-����ܩ\n_'Y�A�"�ݙW��C��)N�k'�޺��^�4�¡�Q\����3����d�(�^��Lv0�����5�����f���;D����I��)cɈ�X�:C��e��C��g��:�7�e��Y�谲�A ��W�TP�Ы.N50��5ՇrX4�=H=�fӻ#J�Ud+�����Cb�����������BZQ��zȂ)i�h�[q���m�c@ �����$
*m��t��	_���l�0��(,�J��G���	���fty_��JE�NLXAG��ۙ�8 ��K��]/$�.e��rY�)�oÝ!�2ل/5�O�؛./�.�0���	>���vfh[�R�h�i7Df�!�8ߐ.�^��
k{<}��)�s�y�m�%˱O��K�m���u�K���h��j�rk�aC�!>.�����@ٙ���}��U����\����^����V�a�)s	�"��h���F_�����}��hZ�C
1J��dܾK1�����i���vC6�/�D�=bd�Kt���Ď+&gN ���kʾ|�=�?m	#�R˼��X�c�����Os��-v��m�vth�y���rS,b�M��]��Ei�z�=�k�;8�\���Vt�����r�"P+y7���6UGaf�%C�%I�z�������tBaЙ�,���� ��dIj,2l����`��|���:�;��l2*���@	�{��:�ᆡC`��u�O�V�ܑ66YI7l6�����.��q�F��@/ۇփ��b�1Y��D�IʴI�#Шea�n�]�g(D�;�ǯwR�'J�r���S�E��(�oE�8o�U��DM�䯤L1�y^�|������#��ǀR��#
�8�U+�mVh�N�P�w�� ��#����+֟�R��oP��p=�� =�.��Ø��l���/�[���{�o<e�jr�l���D2l���
��S`A?���$�;��뱙a�:�~Y��}
�Z_���}^��?C�A�s��0#:�-��v�o��]o�vS�]'.��7�5�]�.6y��We����%���&��Dv=Nԃn/��6�H����C�g�=���oS�ɸ�K�ES�1�wVp5�d�p�1���1�K���Hk S�Y���{KXf�s��OA��e�p't`4C�����,$M5<nD �ې�%*(��0���"��e���W�]͗E�MM+�TywY����:�K��P���r��N3�E��v,�"�Pb5��_ *��"T\�0iYl��=M������Y�zˊ�����rlK���i��}g�	e{�ð�\�J��_񏼙���0�#Gv�4-�o��b�ȒPP�b��i֪�0��[�mn�nwº�!Ɍ�Ћ�7x
%F%	_&i��
���+&6�����G\����,˙"|赿�y�!��KU�������� ƑB�B��(2��y����f:�*_@�v�������w�Ҥ8D�R�@���b���ќNr�%얉V�M�	�z�e�Vv�{�����j��ɿ��R�l�,��Ń&�i���+�`�j���ń���%=��ⱞ�; �<����
A�������bk$���,a�~6�eG
�+��w&�x	<��j�[0�j���d�+�K�FKz�f�"%*#�L�i<A����,HF�5��"��1l4*>�)��T�9gV1K�6>��^R[�+����]�����M�i|}�&pKK��~WC��`o�(
�^��z[;�f�KM�J��1���ŏݑhʿ�����e�ELS��{[�}�{�"X�W_ʊ������A��ǣ���/�?A����#B����J��榪g���@�>��OfIq��Ȇe���G�� @�s7{�W��q2;w�K�uXgG�'Iw�:�o���8�����Yx�>_ÑTU0�%�����	�HD�v���L]Ϭ��?n}q{;M��rksf�� �1ED�.��/M2�qF�LM�b�<���zk�C({Fn\i�Ph��w���;��~����LC��|��0��V���M���@W��g�q4g�ϝ"��!Wy�]]U��l��*���89Z�Z�QbYi�����_8	���6�C����Ӑ��3~�4Dn��Tϓ�=+?���c��[?>8�tL����A�"�	��Tr�}�j�EG��G���"/��^Ux��;��O����t`MƔ���)���w>H7Rؓ����X&��zL��V��@�������Ü���	<v�,BHl�I�Cp�|��,�?�s��=�����z{5�Y���I
����K:*�mN��D��~2���T�"�و�G|���Y��N۵#���Te"S0��xq��*��ț��3m'qoZ�N2P!Y��&d,�УW��d?���T��?�D��ki�d�>����"4~�5?s)�NT���ܡ�]����B�k��+:f��}b4�X�����`�8�Q:;��l禷)B�;�
p#��Vd���r
)q�T�^0�����S	��F�ҼFn�Ӹ��{T�A��Q:<R��9�K����4�/qvX�x �1s˒f�䶪L�a��]��npP��L��2�oH��3[���-	E�@�J~FI��hQ�{w
����
���1�P_8;O��?f����+�T� O�Ja�	%o�oPZ���B����}$
X��3�X�#��M�¦�A!�hd�G�:VQZ]�D��{��xMg���h��>d��;��>����p�/�Q�d�o<�����F��#Q��,o��F�
n7�~C�>��Ga�M�-�W���D�؆1�92o�HFX3���{��_#��@A7�cc�y�Q	����$�?��_b�:b��`&Q=�b%�ȉ�7��A��:׎�R} �Ų��7XXW��'z㙷T�vF���O�ޱg����	�c�����2?U��<��3���)X���OD�Hg+�;�$`�y�*L�Q�/�Vrd&���&ø<�I�b��Y//׵�8E3��h71&,ސ9.���3U���O�!��*L���2��]f�LyӞ��������������p/��f_R���zY��i�;�pw��-�{��b?1��������\�H��.#�C7�R�l���(�y��A��G�J
�-�!H�g��bu��?��͛���p�)t��ê��!1�'�9�o���Z�$����'���%�{�:�?6�4�\�v�'�~	�g���7���$��{9F*�m�.�v�~�kj�i����z��@��}��eJƬ�:�����E���~"s&͟"kپ�l�r��_Z��7��jȅß]L�����m�����Bhp�sK���O�^���	�g�������!��܍�&��Äd��S֎�\�Ƭβ�t�)���m��}�Z��tW��H��w�s��W�˖ǌ����툁2��+�-��9Pi�_Ә��yy$���Bf@<;���<�Y�&��G��]R����8����͎�T��InO9�v|�ʼ��5:�QY�+�P�*M]p_^-ǨVN/�4#���k'�ȴ�o�F}9�@��P�T8;����0JE��ȉ@��"�
����zw�FXeՄ{[�P����:UPs6=������+-Z!�w�$���g:�s���%�3�x��'-C{���>>�u��c����a�j#"����bH(Wh]�N<����M��b��=OcX���URn5|#>�����˂c�n�D@Bh������܉�.)�g4I�^ź=�qV[����V�܃��7�@�R%b�@[_�dͧq.؇�	y���?:'�q����`��_ aG���)r� �tx]T��#�m�q��A2������@1!m0�'Z	�((C�f��d�vtZ����K�unʭ���� lH�-�9A�|���G����;�谅*l��q�˜�l1�;���Vd�&�f��L��t��X)�(70��(��O��t �c��!����Q�4:�_)YR̠������.�7ؔ��jG/�G�#��D�gkIM�E@z�z��mu>��	�{^lZ,u�l	51��Ξ�.]��j����/
5���k��1��+K�N������wM�w�}C�I0�Vi���n�l�4����o<rv\��eaZM*Z9��RF�5�lS�N��(�>�ܪ�J��t|��7(����W���o�D��r���}\M$���^�W�d�����	r[��X�<���!n��2<q�'��`a���̀iifw]��/�0��+#��� �&�w���-��Et_J�B�|����Z��Ni��>TN��%��� l�w����8:-D��o�$�2,�C^�S[[�~������)su/Y��U�QsqY} Ւ�`�bQ
������X�r4˸Br���nwc&m���Q�{���}U�\�5��-����z��X�P�Vo�yeKL틷Z���|q����į�{_b��i��*S��"�%����l�j�Xo+�e�[Ul���7�T�A4KX`��*�7~c�a��������ص͏�%UBD M�O8N�Kn�}�{��M�LV>��	d��vZů�-�����dk��p���p��Q�?q��㒭L+�vS� �R��g����C:'D��V+�!��
#��o��#�"���c����:�f�����{!l	%Aa��8^�{��}t`E3W@\%8l���Ե;?m%����SyG�+�Rp�c��B�Ĥ&�wyoGh�e���f��[>�p����%o!��a�s4y.��d�=o�A�����҆W~�6^���<mV�;fR��UhfK�l7����f+���_�	 "�yZ$�Տ��3z.z\���X$�������>8Fv������{c:7Gke�vk�<_006�oU�ǌ��WXX᫯����MҬH�8P N]�9�&��� � �Be�h�����{�B������t,?}Ji�n(gղj�Ć8;���eW�f� e�"�d��2��+;v͸�3&���+O9���G:�oR�vB��g+Sszh�eT�2r_��z��z'��5�]~+mq�7���������&ccC�����25�;̮g�#��X�s���׼�o@i)��8��˸�{����"WK��ZE���^f����!I�F�07c'�&dL���ȣq��i�:�zp-�?�ӫ'�uc.(�V���7�)E�$�/�2��^�!2�"��R�;�|�Ee�M�dʝ��d/"�L�Z5�4������Xظ���v�-�i}�7:Q�g��z"-��)�&r�p��1�N��4*�8���>�! peVY����J8��q�<l�;�nQ��'�0^/���{��fu�����t����Wnp���z��v�ta~�Kn��c��j�s� �|�G������> �jr�-�ˇ����n�!�Ȁ���F�������lJVA9۴�h�|Y�м�3�v�k/��*�rȽ_c�����=vO���VwB�c �t)��Z��z���^��,���_�d���H�o���AE�s�������p�͓�gd�(#���h��+n�"�xw�|O����}��<�_��d�)����Q��t�\&(�(�� 7�� ʀ����s�|�B��?:�V��Æ�s$+�w�oUsրe�ٗ�D�֐���?��S���#���2����O��5T����[;Q;H�`�ˇ��ܽ'y�a��c�����s���j��}���#˓�����GCl�ɲ��'=Ѡ����^��i����`*"��ڀ�Z����1�-�֩��O������z���EQ�꧎w:�*���zD�Gd�`�<��Lf)yyk$9���MY�3m��+�ҹ�����=?��Z�9�Lu2שrFe�V9�W�"�?�XN�h�M�p�~�ҩ)�<��CKXT�I�h�(+��Di��i9��WQ����� �5���E�?��>"�_��;9*��'p3�i�rg��5��^H�:A�Ϧ��aʶ0|jV�4ä�
a"�؜��а�y�m3�D{&����i��`
l��,�5\����`c�p
�H���)FB�rO����mN����2֧p.�Q�����	�R��M�^��w��ib��>O��~�hKF:7��C�����o�*�/�*jU�8��>{�;k�fi�٣ ͥ��m87g^jM���x`|��+���|X�^)����S�T��O�qĂ�Xx2�݀��u��ӊ6�xߤ��J�E�ЃY��f02��d��20�G0�A�}��}�J�S,w��Ƒv\�%͇��(���1������0�o�R@a=-X��(��S��s��u>\�~/�o-*�'ewzy��	|�%Ǧ1d�z�������Ǚ�j��?�mӨO]Nd����J��e�CW+�D�u'���o�Tc�`}�e�&ME��N�|P}siG/]�ԇ�Y��O�� F��=�����\��7ew��A72�&�մ�6�6C�J��r�$���]���zI/N:l�T/�X�v�1y9'K�=Rt�����-Oe2�� ��z�Y��"��4�����X���,��7qͺo�����G������gBJ� �Ѥ�{Ǯ�es4�7cԕ&�k����w��BG�����,]#������V�}S�T<��y�5܏�	G8�7_2=%q�&�}ì��.��Bd�U��&mt���6�#l��C�����C`�3��R@���R�zE�S�N{�����z?���R�a-cx�+W��4섁c�+7r�?Ǡl:��/:/�V5y�z(%m�6F)D�Cӛ����!h%�ta�UM�H�RzR*[m���: � �h���A%�+��H�����2X���\��[iT��V?�f�Tƣ&�e�Ȑh��N�Wx�k㲄���-��^!>�\n��m,Œp��YF� jd,C)��c���R�w��&S0R������#MG���FmqŰ��ق�z �l��/����%}�& n����ɯ�E�$jW�Dش/9	������byc���8u[���;�\O�,�ą�݃�|�B^ɷ������d{�>˰j�ٲ�M�2�$}]x-����L9W��G3)�	=X�(����E!@��[�^=p�O�r��+�#Y���C���IW��k8��V���t��c�|,Y��`.��Q�@X�H�p��ѐ�(�a��_D�c�Ǿ��pl��=�"@�}"~����d0Tg�ӊ�S@�F���C�	$��j��lK���f�)�Kߋ� �·�{�S�Z��b���kHj�8T$> 6����N\z&�E��"ś�^�F$M~ۑ�G�y��W�0I�Z�@�@���w�OU��Z��՛/�,㢢��/iUV��R���/���i����F)V�^���\�ڻ,z#	�����l��C�#K����O|0����[57jj�h�->���U�a��{[��hsT�� �ː>Q����u|�1�䯡��3���co�E{G��fI����d`��Tf(bM8� �]�׮v��O3�5�;@�F� R�	�e�*�kVݺ���79��"������n5�ԓ�e�q šzϓ���i+#���%{�!2>{W1kl��D���2�Byk� <S�@�m�-���>�k�.3+�*�@S�-��b�|�
g�Z�^f�  
9���=��x)�^.̆o��"%!u��E�7�W|&�{	(�3������ȫ��UPF�����o�ர;qԒ�������:zd�q�{Kkv���Fya%ڶO�F��V�٩��v������-u��H�"��Y+v��]� ��9J�.}f' S�'p��ӜUp@��v,�8�JI@h�g��?��s� ���� �GX�m���W^���De��<�{�� ?�b���#��GkO��6R�Y�ge&9��,�����h�	�Y(�
m�@�)�1n�/��j�繮����͌�C��� q�1`Z�Cp�z`�p,Ƚ��L����ZQ��F�UZ��v,�-�̓(�BF�Y��Omy�3���b Ǡ���4ۺL�v�s���P�dى�ynXc3}���ֱ�*�M~�}H�
���>�$��r�0�?�.�[)���^> 8�a��ڶ��~z�nxF���:�C�
�u��[�xº�?2�o�r���:!h�<���-��1WK�H�Aao!��˭@ݻ>�9�IR�V9���3����/����	J�v��>��e���M/Ԩ	�vuq�u��%靖sm���%��,��V�210{Zq�qD����h�\`y���/`.ö���~8��~'�B���rZ	x�^t�~w�+��0I�"��sV�@��5�>�bxof���cH8R'kp�lG�؃'FeĞv�u[J��%��q =fU՗� �}������y=��➏���:���i�bh;�9��s�¼��p�͠0H�x��A:��W�%J�O^ӌi4\�M���$���ذtf.a�6@�/���s��=�D�1 Ju�������m$�}ƒ%���d\��Td���?�(���MA���-��yP��p����)���:,2z�-6zU�5�b�oS���-��'O��oxg6H��t����^����Dʼu��l����k2liw9~xLM�U?�Ѐ�ޛ�'�`��ru�F�8��-��n�����|�أ@/��;�i��
vi�����'qgj��,T��3.4݅U����`V�-�æ��̄4��y#�8�d��#>o�w�si�=�O��l�pA}��Y�����)�CƗ����|t6��զT� �#��5(!���sFq7BQ�����\�H������N�����n��"s���gʢ.�N��wW��W��Ej/fo��K��]����4����VhbC�Oh����&}/�Γu9����b��HsL��1U������3La�=�#���[gWKz���JA�h��%�avԌW#��y��2Ke�u�٬�q�Kt�F��G���>8P�<��$ޔ��͉I$i�]i]��/걘�Q����r�p�J�֯�*,��Ҽy�F6�����1!\�=`���,�j ��rZ%�T��Q��:��x�b�-"����լ�O(�~�.�H����m��N1T�,�*@������خ���g���)� �e=�mB�=2T�$��N̠�|z� ����!�0�;I���²��~�ɻ������GFMH@87}ʩ�uiw�;P.m���c����<�l[bw�uc����H�����6o4H'���d�� σ����8��쟉4�����w4z���P�W�X�������cg�3DD�LX5����/ɠ����f�p�чu+-Wb�Uu_-�8|%��
�F��D�Sy�o�:�kz��4�3�?Bb#�g*�#���%��8yy)�e�5��"0���,I�0��3jG��79���
gy>�5�О�?��9�` |���=r��ӽ�1dp�K�/&|."g���T�����$�\�����#!&{Ҧ�trűn���u?O�e�h���~�wK `ذycB3|iV�a�f#�X��J,?S	�;M����\åK��7�g�3&(�x�N��ڇf��P��7�����:ߌX$Ҹ*�\̇[�����g�7��|%3�"�y����=LFIz[c2�gSS��-p蔔m�6�b 3���>���� �������X�#G4R鯀�.�R���җ��9?3�u�.ҋ�� �ff��y0au��Ԇ�����$��Ey�5�Ʉ�Kp>T�;��p-W4.�A��Z�	��!=�����h�`���[Ϊa�2B��W9"�"Gl�YJ�QT�}������I?�L��N�� �Ga��Ƞ���<���1���%J�驭!(���L3��
��i�?�YZ0r�f�?�֯�
��7���`U�V*�f�0-m��3�t��ƵY4�37YՇ5�Ν��\C/�w�%C�ěV�v��4���U�v��A��t1�D����P�jfƊ|�j���v~g�/nO���V�L�Q��zkτ�ܭ�!(S|�z��*
����l�D��YXO� �Z����V�n7\񾷥���0���L���ӏ�~�nSB�t��=#^^�Խ��z��b#>Z���} j�{�R,���G!	��B�z�z%�@���^pZz ��"H����_�Fw�lk�_&n6��.���S,��j�oI�?�tf�b]_������:<TX���,(��j&��t�^�p}@�%��'D���ݷ�Pg�P_�A����Fm.+���(�1�B3�+�zȿ���uL�E�$���������i}C"'a��n,6цv+^�<��B�x�3��8dyP��������e��瞭�7)�����{�I�y��T0����H=譣`4P��+���~�2@�]��x���5)�� T���֮7���O�);h����kˤa������B�K(Q/���ePX�A@׏���������P��+M�-�`6<�GF"_Y�$�(*2�����T�J˅��kĞիSTދϿ���nX�cmvՐ(�G�#P�%���3DeЇ�	x�����x�K 1G=�%P��R=���������#�z��2j�k�~4�
Ih[9i�5~aꕋA�f�t���B*���H�/�vZ@��YbѬ�B��|����
�����G�lg�mܠ�S7{��"��a�ˋ	��
Fm���&�i�2I[L�e�<��6TP2��{K4j�A�˴im�˫o+^�sFk��,�9�	H~{�B�����T5qűU&9�����-B��bOm?�������B��ʽ��ىi�꿇��IzN��E��+���u�~w�k+� ����[�#G(�Ն��o����X_rZ�
S�͛�5�?~�[�:���K2����H�`��2`���q2��=��<k\s�yݬr�n�K(��Ъ>o��S���c�1�(��&w�����R�ц�6�\�b�4LL�iZ���5��h��K��⭄*�5l���֠ �g �C�.#H�z�望E(�����^���ޒ����x�d�{U<��ͽ���m>5���x`���F:?�����ѝ�����VZ��@	V�<�#�\��=�_-�R�`��D%k�^�������"�SC檆A>"O��`�岵�N��	�$rJ���j77�Ģ���e@1P�[�����E����r��On�ɻ�i�\O,@L$i�?b���,�� �Ul��Ό�/��`���k����E?U��=C�._,���VE��@m��	���E}�����FO�>�C@̑�je�R����rA�s��w�Qp�T�|Ζ�W1����n�����d��ž��j�K`8���G$��9����V�E+���4OT#uml��P$�e㎙sv+�"�i�py�?v3������D�~�m[�S���K�}��Ig�6g��7��B�\�߳�]��:�9�*�En.7S|����c���i�	�-vp��L��Lj R�W�%0�ԣ�16�ߡ���E/�(��
.*.��PD��7���wP+MS�l�<���U��-:��ûBz%����̏[���o�O�<�,�N.)C/��.1��2��E�N�	�6Pΐ�����F��bLg�}���pm���,2�	�%ny����\+�+D2�|�8`�I;���n*�fݍ^@����2�*qO�H�N�L���]��wR��4 �ÖF_n��X�Wڎ�����Uz#=���:��2��`H��͘����a�b�4C�T�d���U���k�æf�6����3�٢f� �:M��iPH��T�t�_V��D9�j^:য�VÄ�A0��ZZ�&��}C۱������r��#e�C��m4r�i�Mf��.~׻E=�[��m�O=Z%rgK���k��*dK�jX�c>.�� ^䥯�a����UF%�K2��	k3;���Qy�_��;�|��|�~+�~�}Ƚ��f�O�҄�'$�Be���j���t������0��&_]�Ee�L���O9�~xM�/3��t����?��v��qe��EQ��*|��j�K�{K��f�s���o��� OC�c>�!��:@�]����mlP�2������U�*���*n7)�R���=�Զ��;�`趍
V��^��d��?]��?������J�WH[�����~��(��A�y���ni��ʎG)�<��LRNx.P,���D3��/��b����'?&���ۂ��63]�H��㔟"�0�&S���"��$ء��-�&�@�I��H@�H�Α�քe�$Mbv�<�Lc
��n��vʓ}mX����%3�&�|)mSa+f���_��.!ʂ�:<)�,��5�V��!�d�����.����j�n�$�d8�F�HU�|ۃ�ء�s��7�u!���"���n�v�w�(̼��;#�7��pm�iG�cHKS������r�[�Ƹ^���۵��NO\2��m��X���5�(���{nT���ʂe��nW�'��-c���z��Q�ࠫ���/k�������H�e�f�;��43~�`�u������T֟:*�m5b)�ۻǄ�g6�Jᙾw		ʮ��@;:Ȁ V]�3��Ff��������	��@�g���8���V�Z �{;�[�B��.|�Ѵ�3��T�C���&���^| tCr�֥@�4�@<�a$��=��"��Zz:�J�qB��^������.��z@�Pv���[�&��0��ʠ��2j�Y`]����sf�1��F�������:7 c�o|��S��������"��2zO����H�B�)<c�9* �E&�!��x��Ck�ktJ&�����*.��C��� T�)/�S�ӗ�V�&ԕ��yw�_��*�.��:6~���X#3��K���1�`��3$+UJ 2j?�_�uYgj ���MA=DI1e���√�� P�u�H����5E�%���s��U^��z����]���p�m1�Z�Hl�o0�C�ct9#��<�Q2����B�8:�(�؊�bf�[$U,��k��Ncv,��5U�������;���F�ߦ�
���W���Y^7#��	kZ/��<CE?yqQq)�����uyv�4�D��H��k5L)�P@��"�����2�%8�����������y\�U��R�����z�X���5~��Tб�}�=��=+x@�ʐЯ�+]�+��`?̛zJ5yx�&Q�'{�H'�~bPj|��¾��q=�kDh��%g0: WY��|�Ӆ������$�^
c���Q����}��խ��P
b�7��IVH��H2��z�BuGv�BP16�pUӡ_~����X�$���h��7���nu�����J�l���G��O�Ë��D�K;��NO9p����4��l�΄	u$���'����R�f�(�w��*$�� X�K�Ւ��ګ�8�}7�@���Iǵ��YBFz��	�i�8s�r���y %�k�3�"�A�?�q��ݴVD�=¦�P���2��(5��A�-�P���K��U�澳����8��>`�F��������\`�#c��Ƽ1}Kb������p���\�Q��nb#�����	멼77���PULlZ�&cS��"M�#�G������e�d���fM�ś��!�E�\7#�}C+�#���d�]��T�O�B�>̼_�����8��b��(��������tw�N�n��L-�0���;�����)B�ab���ۢW�2SB���$���)k֣��&[jhQ��uf+2G�[��Ѱ�b����S���,f�j�)��I&�
��gk����P#