��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b�����CK��P�哳|�x����`v��&��af����$��u��g	֢;y���0����Ϳ�&;%g�ޏ�l@�
��N��B$��G?���yf��H�s�hVi���h8)������� ��Ծ�V4[AWc�a�w��2B���-lp�զ���{ck^E���ƒ��2<���8w��W��c��T|���]a��NK�� h{Z�	$0���Im]��2��N$��=�T�����U��ϚvpbD�/=��</.u������������d�����] ���L�p~���RQ梲��C����C���ΰdUT�o�9�XF��K��v޼���X2�?��\G_-�6��`�a��!��Q��IO��CQ��A��	~����$6�I>A	���*l'�1Vw�n�i9�����hz�Q��לd���왎m���q1��t� ���D������\�܆��`���|���)M��A	d�t4�/�˝taP@���V%5�S�����6��FpP��h�u�lt�yBO�k�s�J�qS�L졼��<Z����:�ъ��R�d<dݾt�Ăp>#ļ.�h���Vg�H�_@��!"V�X�5�b�X�)�����Z��ԫKR`�J�si�i��`<�Q
�`�]ݔ�����2m잶z'<�E�Y;��(`T�A�PHOt M�,�tc	�|B�;M����H"i�8��D�,@v|EM���[�3=�B�=?_�w��[�`�~$i��z��2B�+H�&��?���ǉ�3�	yo�����`�6�-���"���D��B��C��\����r�%gc���q��I��M]@�-�@����[w��^ٖ����NbM�	sK/4��v���b������yLf�D�Ri��7pj �-�n]ŋ���Ns�4�JTK��E��r�Psml�����}��i0b�r�9�B�� ;>��z���(������;0��,��ɓ]��e��� ��æX��đ�Uۙ2d$�����.��3�WX�OK<]����WOC�7���P�e�-��������$ɼDO�*���Q4��Ae�ߧ�%b(��Sy����	���yǅl%_X�[\D�2�~���£��'X��;��J���!o4�b���H���Y�:����^����$����m�{xh��Ц�ړ�"��`�� ���:~8$���&�2������͘B���k7h�ق_ Њ���`)�qU0�Z��UC,P?���w}�H-.�O���GB��^����1w��?�>�s�I{��w��W9�R���ب0v\1 ���%���eb�&��޵��v�z��Z{����i����.�L03J�="
sz���Dx�߻�>����u�HpF��#ɷ����/�Ѱ��]`�6h�f�[|�����t�`ơ�]C
��MDs�h�6�и_s�g�}����.��f�Z���QE�Y*@�%��2l�����o\� 	f���T��uB�?G���f8���� ����gq%3c򔨘���\����O���4�zO�e��RE�?�3y]����m��	�yÐ�4�-:f:Dp<q�:#[��W{H'���	��'�Q����+��Cx������W�����:��F�id8����O�v�_��Vg���Cl�2��& ��U�h��JSUK�]��a�y���y:5���0�� ���m�5���Q��.�1���*�V��X/EЗ�z��w�)~�H��փ�-ϕ���*i�M��x�x�X�'h�Xn�	w$�ٲ��}�]���YC��Z̕����"��N4����B4�G��iʥ��T ��绱�g?�����{{�=S�����u����{�p(!oq�T:�'������_<��{�8DG��nQ���\��x�d�(ZG�j�:)��� �S��YT�-���������7m��Cexp`isX���h?��d�x�97�*O�|嘻�{R�;�y?��_>��Gu��X�T�6dr �L�x�Eaz�Gq����u]=[N�#�G�&tlƛ8��v�P
*`5N��?�p�'R;7�:ʾL>��t2H�v����>T���3�j����ی!�>gyxG�D���T��_}*�8X�*b�Pf�����&D}���^Q�IOZ��'b|,.1/�T+ld�1�Kp�E��)�(D�C *��t��yE�@���A�-�TֱwF&Q�2�$�nNǌO�t!�ײ��L,��C���j�M7��C������Lv��_���mÁ>���쉱E���(��9LD��6h<g���׻Υ6db����ؖ��'h�@Fpw	��,���{m�j�6GI#1��ڌI��&�Y/�/����ާ�ҙσUUC�3�	QU-^T��B��L����>ޤܳ�٠�\��bL`�Y��Y�N�hb� VE�-���u�9�EE?�T�R����5e�Jǀ�T�Z��f��_��i�!��u0��H��o��ua2\�Tv8���2
7mŭߍ�.��ڂ]�͞�r�+~��v�@Z	��'���OL�8�/�d�ܫ�f �P�7Qa?)�9�v��]GD�EPJ4��
w�����|9���G �K@��1�b,cǢ�
�������J�/���z:�(��ԃ��^��V�Q���v��7P��'����ZF������}�P��!�"�X��\$��:��'n����i��=���As����b!n���#կ��&�8ްR�ps8'�a�,`�Ź��Z�(�R,�e�4<�O�sAߔ�O�9���6f`�R�a��u#��*�%C��֭��������R���٬���F��c�Q���ʪ����3$�uggZ�\:��#8�f���y#�T�G֣]:�Q,�fO:�#a����Tה����-�����~\��E@3=��8b�b���T�;�|ܢ*�$������~�Rv�:Fi6�;�����4)�*İ�r+ђ�L�W���� �qo�S9�:9IY��\Ib�D�Vn�N��E@�>S�M#�2(X�Jْ��I���n�6��3<�鐞����a��SX�����`� ƹ:�̅6h��7!�GH-��z�� ��Ek����j�������S܎FI~��m�,��_rh��Z$��@1%M�O���4�`!��ǋΑ�`����MAS�����?߈>��*�;�n�7�^�U �.�����j,��iI(\ ���V��SEw�)p�¢�M����9ܓ�kaO\߁G�m���tg,�.zG�Y��	�˿���g�B���T�X���������L����)0&W������)��"��6TO��ĸ���%2�����Y)cx��n\���A�r�ʌď���m8?[}�0��J�Y�r^0c�ߜb��E��������F�]V>�������4%�q�m͹��󇆜/\�ZC�\�?<ײP��� i�h�i�H#\��~�|`��YGfrג���^-�d�W�����ֵ��'���#�Cds^Tb��A������e[d�M�Pj�Y���gAK�I,���Ƭ����4�9N�N���MZ\����q��V�ԩ����Q�U�1�.p\a��o���{JC��>�|+� �yxiv�IعSvTU6CII�q�&)��.����]��>ⶠ*gpF��'��+%�3���Yyf�.E��@B_�d�faG�F���n����F��bYX;��V��4o��6�ź�~آ��(��w�Be�z��ͅ��L���@�=x�%0�aV	<B������`~��$��D��ki_;U,B�d���v	�nCpXyC��n�Y�d+�۷7s��t(�4nȫ��_�pۉА���݊r!^K�(Ex�����:3q���$�0[����gm�^Xj�G�}m۞�-�-����s�,
v$`�A���0a)��,����-Ā�xu Ĕj��
��[TE�H�/$��a5i�����Hg���a"�d�y���׹w�Y�>�=�GBtD��
�<�$�mR��F�[��5��,G��2Ӝm�k�yl_�V�+���^����cQ�m�FK�����0x�9�5>��G�!df �+�tN�t����eg� ���r�"�c'�G�+��iZ�@"ϔ>�v�8X�X䂵k88���'k�&��[�V=�I����@�7��D����0�t� �BT�)���x�-I��P)rd}7�@ �a�����,���R��p%)�����N&Ⱥ�nim�b��tװiM�O�D`U7[i�y��)ۿ�2��T�R�hQ����'ԮG`ߑ�	�8xZ�Mܬ9����������Y硊�i�S��Iӧ��(	�-Qߍ�E 8� �=dJٽ`x�(���l'�qn����
U�P����$>���i�<;[F�j�7�X��i��>M�ש��w��q�-�F^=�zC��G��>rS��jϘj �~����b@qً�|������Ԁ�B�r��m۶ޞF_�ނ4���dڪ�������ѻǙ~�,�zټ����H�H�lF'U=�#���/0�T}ǻ�,÷?�4h�{��+���q}+39�B���#�6��D�����S��B\���C���lG��K��8~~sN� �7:�c.m6`�b0�A�J.�Q���2��#���_f�i/}�x��|��s��w�".���O�?ʣ|����s��;�０
�n� w�E18����Zz�K�0H� pqK��d�.\��|���h+E���V��F��O$�8�!{�����UeO�VLo(fg�o���~�����W�M�i̗D�۩�Å��
�_6^gB�,r�ļ��J±�9 ��-��3�s�r4�Z��N�v,Zdm�5��>�eiw�/r���R��3K_��ao	�X��B�����~�$\�wx�� .]w��F��xo�~��������8�6u+/tw����#&�ۡ�	�y�Ν%PUru+��d�1h]숇�΋r���%'(��i�����+:��Ņ�}��=E5�B�F�
AŅ�*���2ۺG]����n�%ƅOVie�{
�,SX�;&�Dǣ��Kt�^��2�O�q��W���x��bx�]q�rY�u��rT�⃂�e�}��o��κ`�k���0���W�o��"���)�wO�Bi2\���!�-�+%� p�ҙ�m����Cƙ"����qW*����h@Xc&n�_�Gt�kX���/�p� �=�JN��D5�}�]�v�%�ΨqYgj�����%t�KW.�5*�R�%ãL/��Z��L~`�x$e�e5�)"L}ᚑ�m�n��ǆ<����m��.r��o\�4���P�R]��Z�����:�j��,�Ҳj�|�g Ӵ����g2]������*k�Ps��,J�@��;wH:���&��H�}:Ѯ^�cv��&k*l�z+k�����P�R\z�zEF�!�K2h����g����-vr|�2m�}��b�*5�=O}�Z5j�z��j�D�+~;eĥ�ToQ�D���7UW������je�{T���~����C�����eM��a�?L�\�����>��f��h@����xlX;��e��$s�(���7��i��t��:�[�d���K{�3����R�w�����D����ota��G9w�S��
IK�B��.1-��<~u1�}���tn����s�	TY\Z���*2��o��-�7�\g�T��~�+1v^�ј���{���w��\|�E��l�f��S_�C�7\:�Ї��ʗai�ժd'�pj����l�z�%z�H䣃��fی�+��h��4?��f~�Ponj��H�d_�����޽�RJjK�L3��TV��CE+)�p���R9��9�;y����h��Δ�2�N�m�%��U��L�.�NR���� �-S�Qo�}@E��φ�,
W�͘7.�ch�pbV��e���F������^��u�߁��C#�O��/��N�T���A�v������~��C;��Y�]�I	�IG�YlA�\�)��>ﺦZcjQ��ىyY�.��NF��zE��Z��%:������=�WY$�p�T��J���:y�>\LB8v� �IWߜ_��}Sh7cTR����S���j�]&[��_�Wjt���Ed�P����.$��8�3"7Rͭ��Q��	�c,(�zE}�g�R�� B���.�Krx5��7t��>P������E�IX�Jc��Xu�+8�@Gɖls�2b�7P(9�͋��F��NJh�gVM̞�Y�U��.��O�9;g����� �TƗv��S�f�Ci�j[�$��GCc(?��WU�ƙN��>�moì��˄}�%Pq�&�E`����a�l��y��N�(s��d��Б�sP̒`vL��)�W��<���끯?�<ռ���kۙ�#�wĚ�qN�W�/.�&�m�i �o�Z��*�ɮ��!zC��(��'z�$!�����KD��ks�C�ؐ��$R5�7jXOe�kr����,Q��;�ɵ�l��-�wI�M��f
(������FM�Ѻ��[���j��?���?�P���9ƣX�P �<c����m�*�P�������Љ�(/�At��j�`dfZ:�BV��w�mRƢ	��)ٷ��������_���f�N쿻e�B�]��v�B���'i���J�."���5],?ӗ�+�hJT ���@$e�d�
6�OX�-��x��J����)R�ԋ$:s�J� �L#�#�rڅ	@�4@FlQL`���!�6l�&�|c���e�!��H��&z��\[>6�@A��'���]���=[�h*��j��s���=�ϛr��Z�$ �W�cy�Zf���7?%����6���/	u�,f�-'嘷?tt�k�!s��g�����.�ȷ�rT+3�~����T��$����ͶL���'��p����v�v�6�qP�
pu�Z�N������7��t4��_C["{��~N�O4>ĭ��K=�z�����h�l���UŞ�n!k!U��X���%qz���{�Q��a*j���+h����+
��ؘB87�2nF$D+����Q! ����/[Gd��4U3��F�8���u�娭p7���*�8MxՏ,I�Ø_)���H٥�ɕ��R^;���C��P���#!9�j�����۬����#��tV���*2 ��~L�����b�g�]��	΃+�w�n�Q�,��	�Ձ�rş�3����C�{M���O���.��o���&^^:f���|s�P'����vm`�E��e��KƴgH%|���&�P�F�E�f�E����&�Y�'���5dA#ae�ň�.޽�S�đ�H��!Đ0�Læ�$���6�&/������ lˠon�h���:�������3pW���#v���%����TJ�p�V�$c�(�'n�!ID	<�F�V2E�Ǥ��NK�������
���(�����ńL���ց��;�cA \QQ	�%�oI�5y�(����a�5��#OT�vN�"�d݃���Xl�}P��;��	'0�EF G�n..>��j4��7�|��<�#�����\	�C�l�cn5��p�]��^�Ni�w��rf��l����?���|1J�������a]�7�8[�`$7��h�ü_����� ���P��rW�|n�4+ub�_�K�(��Ӧ
`5���i&�bb�j|�d,*	���'�3W��ny�5�\bFA�D�:��v���A�vǵ�L�Ȼ��Crmh�b͂����&Z>�c�*��X��ѵl�n٦�E�vT�`��k?E�<��� ja�G��O�
�e+��4/:��Q-?<�[#�
&��Y�{�a��70[H)Y~ H]�akcП���� '4I�������r�"*�`.��bS�$3`��K�j�s�"���8�R�Y3}ڴRa>��Rҝ��5៓�G���A�N������Y��p�HI��Ck���M.�2<$]0�mWw5s��`U�k��͎k��|���u?k���cI� fd
��;�U�R�����}FZ�1��n>�X0����0.�{�u�]��$*�����6���M|`h͆D�*Ik��r.��3���� �L
�)3\Å���!�#�S����y�����k�g7�;���5~����,��2��EMjD��CoO����5��p���
��\�+jh�(Q��=�-?O�=X3L��T��������I��4NFf�Zuؼ@%����"a��B8M��o�O\e+2�R����>�Jz<��K9%�I Ab<F>"�B�ˮCg�gJ�[����;-�$��$z2v;-o�D��>` ��H�|��� ��w3��y�h�V4_��yW�+�k�0T)���w(�����.���F�������E���S��E�p��8j�2:T�ٴ��7vq�����W��~WUXd #��u��3��+�Q�5��؀�J$��ͬ#8΅T>X�k�*�D���N �w�a:�d/�6݄A_
l�({�*4���/�{A�P0Is�"O]s,��-E�pE���FuMi���Qd�ʴ���V�`>�1��o�����"�qx���S'��n��t�6O���DB�a }`B;x��և�п�Y��2�|2����m��7"i/\a�g#\�� �%-6����L���q.�Ÿ�6�҆y��?=�*�6�a��op�X�[���eɆ�eG��)��6���"g[CzM������7�ZY�OaRNx�Ɏ�A}l��HGn2�@Afe�u�;�|D�4vN�g�}Y@�-4��)�Ĩ3�W�De��)���\ם�L�zzy|V��	j9�����mF��?�T'��'k��/�T��Kv#�G1>
���xb�������\,���*�u��V������f�0��VLH��P��D�.v�-��F ߣN׼�}�=�.����GW�����d�PRjb\)/�ƕ��X�c��i���%��Qfw��/G@H��6V^�Z��jb�#�͊	�ݲކ�a��2�������̮�������+!����A&~�c��|w=h�������J�m$���M��j���J�p�#�\�y5�ΦF��k-ٰ΁J���ͮ'���;���&`L�pE	��3�Ӂi4�OGK���IR�m|d�Bǔ�;V�<�5d��~5�u�l�@ik��\�RM�$�\]k��%,6�{�7v�8Hl-������4����n�q���8^����n� ��E��T�r��y>Lm&B��l� �/X
,�!�D���
}�l�Ɗ������I�vl$1�6�/�FrY�s��>�PBd(B$��3F����T>�4N$B���=$C�AWq��!6}%<tZ4��'κ4���=P4��l�������ٌUl���c��?X�؜�g9 ��ț�I��-��ʜy�^��)�y:��M���˸���C���`�jU�L~,6��N��Cw2�(�Ȧ�Â��ם��y�^�ۡ�����a�y�Y`5dn�U8�ߠK�*��+�i����,�v�5���R��e�x���:�\�y�������P�<\��5�w��<ؐRD�H�X�����x��QF����7�� Y��jEDYi,2o�/�H�����F�������#�a����4���ފ"���<�Gݑ����O�d#����*\�#u1#wzcv\�k:#������Gps7�����E���v�x#H�����w��՟#��,��g+/�m��a�Yc�2��Y��ȅ�*j\��3���F|���݉�b q%�A�N�I՟��(�VmB[5��˝������<���p��Iv���B��8�M����.�֟ScT;0{v?&�5�\�'4?>��M=4�����8�!I���������}�R<��4����Yp�C���!���1O�:p�����!P&a�P0�ĺ�SC�2��h��� �/ڿB��k����z��x����G��7�UֳM��?�jy5j�W���4�j��.�G��{��*$�Ԕ�c:%<h�)�mǪ��}@�>s���h��$WZ����P��*��W�}=4�xX�Q%���44
s`�9�(�6�"H�S� @�Z�{�й/6�|{��ZF?��^h��|���?\�aйf�/���YT�)>^<���Ht�V��{v�m�J��s)��G�V���)R
�sr�D�)C>g����W�+3�<�`�Y����HI�.;����Q����i���;�A��IF��*�������LƁ�&A�����Q��L�AX�rI͍-���n{Z7Z ���A���
UX�eH�*>R�pPw��4%�[�������f=������eD���D�X�^�vwI��3J<(~-ux�ѥ߈�^jb }��Њ�W�.&����u����Z6Kq�Z��6�{ãN!ɬ�<��l��+T]û�:e�֤��>��#��g�*)�TM�<B
����I0�d�~�h�9��OS��N����"��Nt��J��9"K삁+"o+�Dw+%��t}�/<�R�f߽���v�5�xr������Sτ�a���nr�#w�d��a	�N{;�w��B���������?I��L��l�^��-��Z�/��c�?�U��'Qs��Ħ;uR0� X�b|��aA���PHttd|�Np�]B��4Zϗ��x�٪�vuV�����i��$7����d�=?� �x��������)�5״c�b�x�����L^�d6`���5�RaC�vd԰�L��G�lk��z!�$lՅ�΁>O��e;jЯ�9�	e�%�A��Bn+��rQ����j�A_@�_!�~J�g�E�z����|�G���`�R,��}S�v���٣��w]�!����o�*|x>m6�\��	��N�Q�P�q�Iϲ��ej��i�F\rݟ��d|z�cJY-�Ͼ��1��ڸ��%�[��ۙ�&ȺP25�L�>�
mO�X޳"1
U�~����Oq������6���=Gޘ��Q���+�'=�FW	l���!�f�����=���+��J	���-���r�:�o�/�6�*�|�v��
�=9J�J3�|�F����:uÝTT��teH�3N^�A�e��p�м��~zS��摘 -�1�\ӊS��0_�;�vF-L0[�׃x7|K{6 �$�&a�q���eh+�&պ/b>�<����R�CI��M=�3'���C2�B�Bp���iM������]�;���d���sT!�����U��W�P6��\	
+L�H�(�XH5�"����VlZ%���y���ֲ��p8�E�B�vx��
���g�����)y	���zq"���Hλ� ���w$�霠�F�$����bz�a6�B-�]�O�1�Rق�F^%~ѳ��!���R�go�d�MS�������	�`����A��}�8Z�����&٬����m��g�W>U}*p�N�O�:z����CS���pc�M��=ibB�L[�
ϷR@����U�|����@SS�u���`�M���U_t���龙���.
@��3$Z�����o��� �{݈��V��;�-��(�Q!x�ˮ�%}?'�����W�-L��5�O�����5ڴ�-��[fӫ�6�@P^��EL�,[�%~ERr6�[����p�?���;���a�����l�d��z�P��"񋤺�U}&�r	��8�{(�n���w�lÞ*�D���><G>��"В�W�N�r��KiȤ�Ѧ%jG�̄�I���D9Wb�(p�B7��xhؽ�7�n #�[T�&�}�T�ڑm��q���2sY�e�Uun����\�+����Y�89xA�a��;�P��g�1yA�a�,�ϪQ�f����Вqx�Q�.)ŒZ\MOw��\&bB���Z_���%tU-�$6�O�@��%3��w���|S��%߸[�B_�[U�A��>�WR�S���Y�^����0�*���>��S�(fp�wI���=�η����bEȂ�T�
8�<�ߝM�pSp��ҋSEZ[1%��ɵt�N��B^�z觰3�_�h_�)hj.~c7�1���<B������z҂�248ռ�,u�u����	�6h��o���F�����(�^����4����kmu�R�B�-�S�YMk!�-F�t���x�H-2�-���ڛc���+ҩ�����pz>����t��5���f7NEE�Q���'|���P�n���ΐidmo����������칅g����]������@YU���K-��V'���U@�4*m�z]un��8�'0fw��r��W�v{�o';���y΋���2�ͤ��~�ǫ�ћ&e9��]Og ^M3����f�t��my��?n�+��;����A5��"b�D�,�� ���� 
�RE�p�=?k8��mC��$l#Q��e��]�'?̤1�"��au�nV)���N�U�T��"b�zJ��'��:������=v��A�:��A���OlȮ�f]x����Z_�T[�/ǽ�4��5�&�ΐ��J[=�D��6XI�Ɖ�dAsԮ�!Z�0;;�PrWF��nT�1D��m�x	�L��8 ����&u�S��k<g������!Yu��fM��5�����/����f[Ĥ���.-I��J�{�lٴun*1��{��3z8]�.���|��� cՍI;��bA�	�]{J�cv�+#���ր�Ac�� ��@3��zTXJ�7H�e�u@W�UK�@���t��x&�q��|����(����(�������>�o�����+?y��	��=� x�ܡIȗ�ԝ��۝,������n�Y%n9�pM�	�!��b��z��ߝU�fo�D^�hˉ6��e���b�Fߗ�O��bm��v:ߵ�Y�J�p9�c��gӎd/"���	`�YR}י/�T���-�bD]�+z:{XN6l�{D%��$�#*�H��x����[$�zݔr�V��F��Θ14]@�P��8:I9�a�s:�CT�9˲��<�'{�eb��Y9��7�C�����o��t/D� d0mc���U�b�\�]�,e�;S�DOG|�Y��rV����� �>�b�.�9���;���c	�?�x+�"�Qw{��o/�).UUv]�*��o�+5"gKL�2�;�R�K`=|�y�%8��m�;&�X��`EJ><93�Sx�z�8��T4\!4;�;�}6�%�Ĺ.j�����+�j�n�碊?������[�T���.GD��p���Œ}��na��-�Ԟb���1�c�eS0�/��I¨,��=f����e��&j86B�T1��x�I�,��l��D�2���3�H���\���@�uw�����6�&Kfd� ��B,Zz<�H�z�ƠIQ)��N�:o^�%8��̽iGr`�n*���G�5��dY�&Ķ�F��;1!��Пޕ�T��;$y�W�4��(�RJ�!��vԖ��B~>_�Ѩ�� k该���&�EDeɛ��45�6`0����:�˅��SM>����ݢ�n���\��!���6cǒS�pp��<�G潟���Q�/[��H-�{bn��9X�_��dsg}=3Z���\`qr�b�.4����4�$�m�4��Ʈt��XnI��*�;cw&�/������}�O	�R��)c��UG�̋ڭR�{��q|[��?c��T��B�;`62�Z<���n҃�����4��J)��|�aK/Eh�hX%"�<��]�^o=f�hK�4[�(bND�z���ϗ�8��
H�s0�k#C����N�0����e���)�,��o%��_�m�}Z�\!�_syS؋ ��\	VU�}e/6b�&!3�VA�{���&�h60�g�靭zi}�ZN��a�͹�vq���0��X�c���G�H�"��x�ЧI��iXx��溉+}�S:�&�q�	��1_T9�[ 膬��l��7��L%JWԏs��:�r�>��F����5'ǃ?*y������>J��&F�̼,����hr�+p0TwS�P���U0g��ҿ��e<�]yD9G�e���#���jeV���G)�����	T\R�,G�K����8G,������z2��w�Zd��Q��4'��Hf���%)�$��,��g�
���aj��G4��w�K��.y���=ļj3�ZS���T_#�}8*�q�{-����>�V�^�/��J���C|V��u?�����Чeq6��c���ŕuO�Q�郤�_�>�S<�mc�S��ʩ�Wݧ�!�F�~Aw<V�[a_x|2�+\��Ļ�KJ�t���ZP���n�����0Ƈ,�_[�r���R��g�/y��]�l��}��d���I�nu����<�N��? RP$c�G�2�^��rOס���B���U�J���B��Q"S�DSf�  �x��JhE]�f�O��MA+�k79gZ,��&�Fa��O���I�2��1��X;�����6�ō��sïzJ�kI���N��N�������!%��t�=�c����*�=��R2�P�IՖK��a9�f��[�B��KY�EN$����X��12�Nԗ�;�H�Õ��0�Q�@������2ϱ�n��<{LF����T.������JP�"�.�S�G��[}��K�����^�b���b ���Ջ�Uf�s/׶����>��ע}�T/u����W#w��w���cU�1� �m{���X�>>ya�Q�8S�vO8[.T$۷������j� Ne��-u������UW��s�}��߶.��Q&��;����#_��۞�����A���#�D9ʙ�8�J<�
��c�V�P�R�����n���n]Ȟ<;��IM�sh�{o��f��}�9a�~�n��OƯ?	�fGz����2����g`u�a��U;h~�.��1h�|y�	�{�N���Tǿ.�U���ھ��(�P>[D�I��%�&�/&0}��]���	�ˇ����i\]�ܙ�KRѱW�<[�A�I��<�ݶ��L��P��ٮS:p�(CU��;{�������_<����%�o��c�p\+m��b?�25l�~KA���X@79_��yD)IS%�v%3��E�Gd;A������h�@�g~]ɒ����D�7q0l�t֕��ЗD�a�4�TCN�l�P3����x�G����R����4��lք�1�J>�:�xp�*7�ZM^�$�k��Z����iҟ��~$��vVS[G���e*m��x8􂋜�F4�ɕ1�,o
�:�m�+I�?��ִ��� �?���i���*?�v&3O�]���Q�,�x�~�_�����B����0 ����>��|Y��,�xC���[4.S�ŻK�C%��b� �s���j;��\���g]�ɍ6X˗�8.���cf-��;_oA���z��~�n��˕��l�H^4qGc��@�&� $65�Rr�Յ�v d7�a'?�R��י�æ��4sGn��n��UQ������eTu����@�4�M���-�Z�>9���c�(��Q �IF�-��:LQ�I؃�a��.'�C���}�	\ ���7���J�6���'��&<b��� ������{���+��p��b���p�N�������X�4������f��F�2y֐ήD���~H_�c������f}��8_^W��v�9�A��v����d�]l�N���k,lјﯠ��r襏�(%�/&:���W�8B�<��ߧ�k�d��ڈ�Ӷq0'u ��q5Tϰ��C�ڽ��nk�2��z�3��VaO�O42{�P��]�{>�kX��6�٢g�Ur���c��T�X�P�l�*�|�iՈ�p�&���@��N�u�J�-da�f�\��Z���w��"���n�4�ڳB�rR4q1�u�ר��X:�R��_ 9(�s�߿�� 
�_V��3��+�o�7�!2�n�es��>��:X�h�'�;�a��JE|E�_	����MI�%2KJ e��tu؃�EQ��<��H��E�k�K}�f�d��aY7� #}���>8d���6<�Z��/��g#�y�-�VV�ұ���l�-��9zm�*�:ďw�q�~�	XVMb���Z��H�bI}�I�q�H�]d��� i�F�#@��ǙD��J�k�Ċ��������O�|�Nq���	C��P�'�UU��r_��΋����2B0���?r �o�h�<et �vXU�;gqf�=��,���� �� ��v�Z�r�("���=~T!%��{�8ad���������*�J:\s��G��k��®��;�jԫ�
��^���gc���"�5P��.���'����wN$?*���  ���yK�U62��Q8A��a\�a���䟵*$ݪ���i��� 23�ְ��愜Ӛ6�H�v�#i��Qjo<B|8�E��	z�X�U