��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�U�����w�7<@e
��*	�E��&c���:�2�fuaM��)8�C�x�j��C��g�+��k�D�FP���]?(������/Ԝ@�s�D�K��Z�dp-5+r����vl�7F!�e)M��Y ���I�)*]�1�<�}ڲ��p��#/�[���a�Ú�;~�#�ʝ"
A >@i+s��E0�kJ�C�L���`A��+�2�s�Fz��k [�����D�9��n�h� �c?��#��#)6q�_��-v*�hE���#/��%a1��}st#�7�>�Ό9�L�<[��f��r��?i����J�� �mǥt�*��[Q�������W��- e�J��7i��n)�dj�F��;��za�ϟ���5t��ޑ*�O��.���g�t��+H�j�.��U����>�z���Āe��}�DUb���} �?�1F.;�*"�+�\�ى/�2z���]DS��f制?�i:y�^"�;��k���U�޾U񩦦��xffG�g���ENո�խjuҸ�fgA� �[inEp��ͬ+_T�~,xl�*�T{)>�֘Ixz�N��:��Mr^�ro��D��<�x�R���e�R�!r��=�:�1b�4:qB��$z+�R7Ҳr9<�N
�jI��\�׳85���|�Ŕr����f���z�}�}Uƪ�&4VDg4{%���߇���ɣ�LE�tku>��So�+��3v�����1�Tj�+)���5���z&u^q}�(�P=J�.��|uL�����V����aj+˰�����A�Q}���l
�cn(�@��X6����/{��IPCѕ?�S|�N��GQ�*�Mּ�HRj�'Y%��o3T��6��Y���o��Tń�D���8OP:���R{yG��H��u�jH�E4���:k2��u�j�,�ohű��V�F,Fڑ����2E;����n�y60�)�i�$;�>��-�l�Zi��9lW=�.��9��W/���WFl������Y���pp�H]
Zd���{���_B���!9���}!voոDӣ��[$W�:��* ��l�K�pGS~b�ֶQw��KLM1v��ǤϴJu^<k�9\��sWPLwi�m,\eC@���Ǝ�*M�S���y)�t�\���]UY���� �����Y�r[�ha��QT��l���a&J��������,�E`[�ʑ����"K4��::g�@U?I�s�Ee\Z��}�7J�ߊT��[g�5�%��k81Hܒ���Ȫq��i��>.,���"�5�FP�4:���nO��}� �I��P��>�<�P��ͨ��[`&!�4���Rt��8[
�,�|l!�8�L�Ϸ��9����a�FY��HOb{sU[.^�x��i,�jq��+�D�Ba�$EL��a�q�X��e�;�[�� �L���n��l鸙�L�̂p��P��!��e|@j���N���ũ���-�:��Wt��{VAp�)d<nI�ENg��r�Ê43)D�C��$��'�=Gb"�`� CK�[}��(��6��|�9���+M\���g�ge�T��XV/-��,%6G<ڱ�˪9�k{< oH}�%F�q����H�q�٫��r���Jz�b@><������/F3r9�q�\�g��f�0���"A���G�`׭$����O�\�G6f��Ɛ�"*�#IU��u��w��Eû?�>*b�,l �N��l��{+s�#`:�.�����ߧ��R;����4�S�^�*F�8�j 灧�^�4����YG�2 �<�{a���LB͑�\�l 7N�%V� �@lk �����Ss�������]8|٨5�1u9�b����do5�<dګX.�v�,�8�k��W?�����:��;���ȭ�����/Wz�
kע:
��PQ�3r9�Y����XU*zq������r�dQ�܋�6���`����ެIM� G����3=��Xɝ.֬�*����ˮ��9U��)�9����O�^�G���#�N�8�e�OY�|"rx��q������$yǁ�h���[(U"tG��0���fn���,��"+��Sq��'��k��͋��ѧ�3����n���%���?>�#5� Z��ޑ�sO��
uֹ�.g@<?2p�����uuxV\M�7�D' ��/'eF�q.t�ƈ1B_O����tYmH���E����$^r�~��!���J��'@;��TlW��̔f5�H�{�`{���H�|QB[E�!t$����)���M��3����6H҇�'S���rQ��dj���6���]k�����YМ��nwR���f.���#��kZAC""͝��ۨ֕�e��0�/���uMv�d�P�C'd��_U��L�X�Ъ{/�o(���Wa���g�<W��ѡ��SR���LZ��Ϭ^�ve)�j��[��?�+�G:k'�3]���nӵ������yç����H��vT�}�	��wn��Pj�a�76�Æ�V4�y�oϕ��Ùe�"L��ݲ�|��ր0F��@ e��is�6.�t��7u�JZܐ�cRåŞ>t� �Kz	\����<�!�0|$Rѣ�Ī��-�~c��u��^c��L޲�8<eZZ)$��eɮ�N�~��A��]��s~�o��OQ^Yc,KV��!#Z�^��*:gdV�����QeKx�92Ҽ��DVؘ{W\j/��I
� ��B6��Z�¬�%/W�>r����7�i�Oԓg��j���\CZS����0���R�ȗ�(�m�		<R=g�q���D�$-�R�/`@���h��B�c��:P�7xY������)�T�_�ɶ9)2���	���-����2F8F�Cz��ҩk��y�\,rޑqܟ�y�ܔ��Q�	����6�4^vDw���6�Ny1���Y"��M��<��X����g�~�g�����;�� ��1
^�!-��>�og�k��h������↜�0�s�ah6W��������lP�#S�U�w��6¬	s-��߸Iat˱G�Z�S+�0ǲG�j��ZDr��(��جּ����s�2
����`�y�'��!�Ë4�ͿL�ol�aU���8K*�e6���׳���������U�L�wˌ��=y� >���+70,QB�8�=��l�/H�;^I^&���H��L�Jo�>�I���>����}��	��"<��Eo�,B���K]�]Ԁ�`_�i����#�w����]l�
�\��$�,��i�z��J�8��3#JY�2Fq'��V�)4R]-BD�p/��/҇ ��{���7�^.�xSSQK�*��N�3�XKA�R@�ȩ�?G�L�55Vg���W�|�k�|t5��F�b��<>�������9��aw=]3代�1�e_�dC�9�%V��#j.�p��~��|��AE���:�o��;���EYL�=�cN}�w�h�R��F��O�@���ѻ*�/n3��U��+Q��*���+c@��A\"�-2��s`YRf�9|-�DLZO� sTg�;�j*#z�����W�sOR>L�Q1|=~�J\�n����jG\�i
)k�Y,�:K��I)Ut;�@Y�U��1E GD,Ws�����?C�\�f�4 IT3��(��Vcg5l��kw�����`�=H{k"�W��i���m�$�hn$��9���<�K��]N����I6&��>�°U�-%I��	�=(2E����(��XpK 40�R�����2�90GF+~A�ߟ$t���}�*V���)��:����*"y��+$�NԬ�&��v	��FF&���S?T�qv�"�@��j���{��K[V��%�>D1+,���*ٱ��_�i�]F!�I�%��?v7R���n[���JyU��%�"y!��������<��8LP�^��P��;���:��أ:�L�p���昳��b{R�@H"^�&}Xt2"��t:��2���V�y�5}7�0��ġY�f�L"������e���)�Cѝ���>�P:���	���7W=�r=��=K��N䪪�&+�����9,��������FP�(�<g_�C��\���J���P�EG~m+�A���9��fxW�y�����`V��Yh�i<|Թ�%�l�h����T#C	A�a ��ʄ~E}UV}�����!K��N��{&�U5b:��k:ʾ�*/� 	c`�z��AB�]�fm ĳ��e��@��xq-�Z��e�n�.(�C�suҝ,�C_e�B�X1ۇ�;�]�������X�}���+���<4�����z��[�g�Z�/�*"������,	��rg�Q#J��� He`y
մ��Y#����h��;8S���	������S=���u[�X�Y��,��1��+�\�q�~"����i�j�*�D�Z�W.�_�,�νCf�.���DqC���!�У�� �R�@�)5M��ZA	����G�f��$�%y[��<�z�����,����]�3Y�~=�"�<l����@-F/�~��Z���=�=�^��k��xA����l����D�(��G'��8t!�%�F^�+Oq;0�\����~���.1dKN��nS�����);%�w����E�Z6�(��2͉ȃl�v<z�`�W�dNe��LP7��)dQ;��ݰ��� �A�~�d(�l܃bU�ƪΓKE�Wރ���.'��t�8]���Y?��-����v���Lǡ�������CxV$n��>Z�"�ը�dc�=A3c�C���,�Bifu	�,j���8�򽜦������:+�ڗ[�gFf�xq���V���o�|>Q��E>��Ŏ��-!�b��|~��o1��@�wL�'yv;�k�A�ڊ����xׅp�8�F�5����$P/��0��R=�[UO|�hv���!�6-�].{�k+�#��KL�?U��=����%����X��c ut�W��{� o��]�?ck�eot��d`�$�/�GhA;Y�!lS�k�󹰒|�7���/ٖ���;�&'��,9@��~�Hw[EL@�1�X�^K����<%�K�;�{sD����	Ögfa5��]v���/?&�������O���l��rٲ|�LȑBv�PK��B��	A����/s]�L��d
m��}H�ل���y!�l���m}-����ݎ0Rb��a�a@���T�H�_#��Dي'�����qN�鍒��Ɉ���� ���H���򋕛��p����׌U�F��ŭ]p�W�fI��P���ʢiⰀ�)B�..mŊ��ɔ!�#X�]��s�d�hd(��g�p)Z����3�AC�5��#t���uH����#}\��ړ\���q(��3l��'K2j5��#� >�59>���7�ʺ�	�'1�q y<�U��O
���~�(�}����-q}!U��a��82�3n<��"&�gp�O��E��a����ze��Pm�u��L#��h�~B�+�4I/����o J��Q4��L7�)����?=����ײ��wE���^�e,����,����|�]��"~}�?'�":y}�C��Atg�A�����m-�5��c[��rp`��2���k��=�൱�w���=�w(b�I�bӳ�vIq�|3�50��FFl��Ey|�ϫ�_�H��Hnۿ�3�p��/hG�nq��wy�jW����c�(�9.�$�~�3�b���*�} �N��[{����ߎ���u��|D.Ӣ�:���C�9�����f����ѫ��V��K(d�p;�Dz+�P�q"�-3&�6�}��2NT�L�q|w`�r*w�9��f?_���k�Pj�1����i���o�^=�{���`j	ȡ�c�����ݱ��?�6����V����@o-=P��N�n�t�{8�t�Ġ�+��'��}RsQ�ث��y�B+��h�ێDF���M���v �i/�[��
���Rz��=�b�g�{�o�Aڡc�m7tY�׿}gyv+l��ǒ��h{�w�����pL��qf�g��@`P�uኢ�w�o>>R��K-��ʝ�A�K0 �[������W�lbRO��\C�G�zx ���%��HN�k�_\R�������+�zoˏ@*zcI�í��[~y��R��v	Lӑo�jz�R0G�	�,uc3�e��_Mn}n7�[K��O��bD��d�����'�g|�YUr��[��Ʒ�B{3�|���[�-W>�ӱ�R��c�Uo[*�Av�z(+©��[0e#���	x6�-�>�޴�i�G���w6�N��Թ��S=���(�R�+�idӀ;�/�:w3i������.�jt����r|�tC�y�x�����`�j��XR���e�t�u��S �����7�W����M�9�VC{W��;qF&��8Ԅ�8��5����j�����p
V�Rb9zp\�7�
�m�?j�v��?R�/�H��uc���ϋ�4����w�!��1� �>�2�i_�#JT_��^[Fr�_$F<��]���Y��xڤ��U�ʭ��J�.�(�s���&A+��jTSX�]s'����aHc�ĕ��HS�ʢ���0�$�x�S)�1հ��b�ǔ�1�䃯��zm�Os�F�!���?��$�]F��)?ж��F@����K,�ܔ��P�)�Û5�é��܉Z�������o5b��Α�Y���%���mE������6q�9H����Y*�N��Q
@������ 7�("��̛FlBtq��]xw�Id�Q�UA.�`�+a��g�6�&��lOq�m�r������!�פ{��>���\i�L��G?�5sc&��mu$=st��G�8�JU�u��U��M�xz
���,��]c{ɮ�X�����˥��\�S�K� �O�ΣN琅����έ�ݙ���:JNuI�=d/��Mfn�� 0�ŗ3,W�sn��	6�.\iow2h� l�MN��	or�[Fԭ<�IG��3>�%�E�*��$-m�B��f���y/G ��LL%�F>gX(�P-�	���!^�s�(D�䡋�(y �NN^�.��IH ��a��\���"�H�h[��ך���t���)\���<�!q�S
�5�.��s���S���<���xYK�&�3hE���~Ư��K�g��;GM��v�k�Qh�r��w�O��$\-D���@��IK�]����RT����R-4���,Ã"�,���*�G�Y�t��u�6Vb�y�x�r� �A��=&5��Q�Ϋ?\l���K�?}�$��Vgd{2������&O��q8h�>B���0�c�:h�t`�&��3oP�X(=R������[h]x��q�+V� ���3��T?��:sA)XEY5v5g)�z�����+�0.�׷&�1A*�>����"�"[���Z���ȳ��K�����-]\"Ԣ��]gH6wdzS�K�m_`<�6����O��Jo����z����8=�E��_-�-�	;� =�t�J!9JEi?N�3^��G��j.^��0g9�Ԇ·5hc���%/��TP#f���������h1� ���~$��)Q�vD>��{x����f/�vP������w�&t�w��jP���:���͆.7S���j-�q�-{`�@Ȍ��Pzd��*pM\��6�:��R8�j�R��K��3��R���3��0k�E	���T>n=�����D�l������+�D��0�z��'l.���9\ʮ�qa��ݮ/�4~�A��mĿ�ԭLLR��\�Gn���0��էvz��2z��hI�O���ݕ��C �����n���B9�H M�(H{�n�Q*����P�S� ����y�}�s��u@l玎%K��rh�豚B���Q廙�I�����/�bA��8��F��]FD�����Ѹ���׹g���F�_��2��A�D���+gޘ� 2
��0�X�u;�>��
�����:A�.�2!�R��9͵`/ܙ��b$(f�1��N0ԢFW�'$L�8�z�Z��jrJ�}4+�2��hԠ7�I�h��t3�{�_\�B`���Q�2(�7��.�i��G~O)G[5�B�3z�&�ŀP����2sF��M]�úB���[��#eHx#+Z��Z�o���^/a;ZL�^�0+�-�����=�xe�{_I�*�RH�Ԥ�壳�(?`7����~�t�c̺!��s7^9�G���͑���+��֣f�5}y+�+3��jy���t�|]"�ûuX~��'�h���\N��i"��e���Whߥ������� {��ّȢ��0$D��؀Z~��vi�?cV>����ͤQ@4{}�D�tPt�UR�2J�]���y�k�����g#`R�hF"l�-1�*+F�e���Bm�vA�&f��Lؘ��5��?��H�\�8��f�պ�k��`%�]k�n�g�R8�k�\�"���L�.�I�IP.�*b��A]�\_�l>���t����=�EBó$�z���~l�*PX�E�W��ۘn�,��n>����[��C5���鼟�9-���ml�i��ދ���0r7Em�0����^�M�x\�׳=<k~�f����׎���;��<-��	��g'D�n����	W���U]T�~��=TS�y=:׫߇[d��y�����͌�N�9�ҫ٘U����jV��K\��H����&�I�6�
��m��Ľ[�lM[��Εx�D؟�
%s�:
����J���ca��j��;9RϬ���ȣ�E��&�KB�m[ϕ���F�#�����c!#]""�EOY���4ۍA<�r
y]�������|?��lF父�K�}Q�X ,�q�_�(9�{�K$#� �;��`���DIp���t��H�;|ԕ=�ֻ���D�����ZN�
dc]�@�����
�X���5s���Jg�RҬ��Ip�`㓛P�$+�0�P��]1��G���Ib�1�!���h��(|��>[:q��P�u���Xw���7����Y4`����~t�@��L|M�3]RA�Y�)�PS���g����(��7�b6�?ޭL:f�k����K
.��d��ڎVu��%l$]���d@��׋�)�-ɵ���>����R��7΋�@��a��(V6�k�wDf�8�?G"����0���x�"Q4CS���@\�\�V��;W�����`'{���ZК��,��q��&Qu�ߨ���k�J��
��u�"ݧ�%/axd���+�βg�&���̔��Z��r�P�~,�Nߏ`쏱`^V��e�n�D{�&c�ơUn�m��k��D�}w�́�7�T�^���PL���0,sGY�'�F�,ޙ�K\��By�YDw�A/�΃��	 ��{��<��Z�T�v���Td��pr�G4�Ɠһ��
�F�P��Bm�%iޚ9?�6հ�I�w�2zt6[��R14��vuq=83��y:��%
�Ҿ<^p���+;�m-�/��0�?z7�u����� �B��ɢ�Px
S ����	�wp�N��ɯ"�2�p�7���vH��P���?��=e�)D�sՁ��%��<bn�N\�����\���|����a89&�0E�Y#~��imp?���߸���^�LٴP*#�qWO��!���Z�����������i�b�w�dʪ���;�.���du�Hye��J�x2�fپ�e7Eֳ�:P� ��-%@A�F��l+ ��)N�e��.&�/������q	�%�l4cvup�_ǸI q�4-'4'����]>H���6#���� �C�3�\�㱫�#��0!�հHq�������yʥ����3��
�3d��Y��%��~ �g��c��v��x�&G�¸`��tp*��w~��� T�ᛂ����-�R\��v��fgW�(�		��9H	�����)� �~u���e�xgT�u���K����6��WbĲ�H�9�)k��ر(�ĸ��+0/L��Bk͛�fXW긨�OaN��u��T:H|հI)OIbeq=�w��2)"�s�`p��_w3�]��[�[�h�a�b�9'cq�ɘ �c[ |70p�����И�+����SW�'�ёNL��,�B�(�jO�BF�#E:M�L�Z��qc�Vf�&�׺���&8h��Z+B�U�d!`���:`�h��K3��!"o��m̌�9��e����й�l�G亀t������M��n��268��@��!@H�;a� g	�#ZH̑ ��р�RPC3E�t�J�6`�q�%�4|�4�G�M�|�.VQT��EPecl���E#�K7�K�t�&��._�Vߪg��ʓ��z���K~��VJ��)���6�^S �6��@�2���~�.˫�ʻ�v�MF�$��-�lx����D̵�w���_S�R]v�}"s���}�2�Y����@��O���~f�S#u��z�W��U���Hcѐ�l&q��M�*�I\\���Y.ʴ>�w~L���1q*.������f[Cf#�u���A �d����P��50��dj<�k�O>}	 (�gm6�B]/��ua��}٫I�]�7�ĥ�z��S�<�����228�-���=�� }摅w�؄]K��M@������<�G�b��s�r��|�CJ:G/}�'y��0�vI�#�V���ݩޅ��S�HٻH�A_����a���7=[W�e���P�5��0�|cd("��*�ZÅT�wC�Y��Y��Ԃ���M/%�e������N����d �Hg�Y(!;�r�|�sA��f#^ޯ�� �>]>6�1C����x���!E(��X��$\��@�H���PG��l'*��H��FAM������y��,���1�B�w��Ĭ�I�:���+��f��+�FFW�Yc!�S�(�SOQ�Ѱ�����V�xl]<�%^R�-��8j��5ۀ6�����F-> ��+eA��l,�~:����Ű	c��p��cDpN���x���F;��V���a���g~�H�6ŉ�N�!��{�֖㕸W���e�B|SO��Ci������,�1�x�d2��ˎ>!��?C҆�2M��ԫc9�{�x�ҦdJQ @����*^ͱ�@ɪ�d�qz�m�,��D�74���L�ro��p�M�|a�T�\S;6k��z%�0qy/�������`:*�c�c�;����ZPZ_�	�&�;8����P�sy�?��g{� rd�f�ʓ=5)1�R���2�P�x��T�Ra%�j�]��Gcr�*�Z_��"lG��9�=�]��2�_HDVҒa��?:�ʋ�c�)�z�-���K�q$�3ďt!��c��'����Ъ��˝�I� ����aEiZm�\d��p��n�s:��<���~�짍��);!�U��pi��e��p��b0q�=^�p�����@K�:a�J}:������%a���s����Iٻ���4sY�'��$uX�"�q��EE�qM�9Q�k`������	n�g���
�b�W�/.6Ī:��Tq�v�]\�pO4��9�KW+��	�SZp����G%ŋ�}6�)V�C�@v�m�J�I.!&�ʯ[/mz��e�zF�$�Q���%���~�	��"K`���E��%ff�r7$���.�=��X�uY��r���5Sc�l�G\+
H�g�R�5�GWN���J���/�[H0I���w��?��?�D�}`�ds}c�H.�/�n/���NxZ�~���v6s��E�S|�1��l�( ��@'jl�A�q�_�b�!Wߦ�o�2���`�6}�&$�a��ޭ7#�Z�g�w��M,b7��x=���U�T��٧���!�M��'5�Y�f��wC:e`����Gb���>߰�H�8�WknP������U"!{q�`��Sσ�W�mT���6���k�a!�
�������p*H�Tfn�����e�{�� ]rW�v�}AN	�,��{3
��Ǝ�T���FZ��u�f�^.���Kf/�g��W}��+�.���L!��-V�-;�A�]e9Y��� ����2�G�`����V8c��s��=�p� ��=O��~��6��D�2�iO�����v2���=��,-�M��s��sܯ+��Y�R��F�H7_��Ӈo>@�� mCimdQ��/l�#���[��h[�h�n22�����h�=�ڐj�h~zƣz�Y�i�Ҭ�L���C�vj��,�4<`�ì$�]LQ�~/TT2�� 4�����n��0��E���}U��yh���*�?��o:Ӕ�ǲ��h�*b~c�/���T+j�Ɋ�F�x�\�]�!iЧ�⸂�KP
G�)^ˉ���T�İ��o��+� �u#VF/�yE��,���y�b��]��f�B^~��9W��81�_H�,��;�o�E�d��sN(�a �B}�n��i}jA��cc��zTfY4��ŀѭ_{ �RcgeĀK4�L �|0�z�&�伢��h�l5 ��{�a��E;B��f������g�����dT2$6��Ä��tnN�
tC�hmb�Ƌ��{"*�9�y����;}j�}�\�̦�`�QL���&�'����7� {c��O��mlLK+EIڱ1Ŧ ĎL9r�0i8�iT@ǆs�-�I�/��81����9s ��ċ���M�o�_����%vE<J�{��a�w�DҊ�s�э���Fdǵ���!��(Y蠟�5��P'�	��}}�tL���}�_&dͨ�Z���w�Xðe��k�s�#j�y+4����Xc��~Qc@�R)�>A��r:hKܴ��W͘�4�,�gʮ��(�8"�/����C�._<�K��cCz��w���χ�z���\�߆��S5����DF���e������X�	��.򧠛(���s���,6^R��Q�Rǥ?@';Yj]��h_��������sS���w5�F��`E(qk�q�!DI�9d`��$"y��y��)~as�����|�pο�����г���Id0�z@��I �����P	�lr�t��_�M���.�UX�0v���!�nUe�	[QR\�`
��� cg��;TZ_�!a�A ����L�Eg)� ��0���gߗ��6x���e�R�v�  Ӟ2_��,�X���7�ç���|RY&�8I�*չ��(%�r@	���Է$�'-�M'ZT8sd9��1N����E�_���U��*���XD-G�ʩ�C�pU�z�g�����*��w���P���&ɕ6t@�Z�5>�"ڛ\<�����0k�~�l���M���ݪy��M�,}Q2�{�j�bv�
��aE�t�ڴz�G��_�U��wR)Q!ރGB�-`K�{U}W�_lw.��&x��	���&rs���k"h�0\4X-'�QÝeLkl�4JGz& �_+ғ �g�v�����qXQb�����Cl��R�l�2p�3���@�B�KQXUu��D�kEnw�*�h$8I����*�G� H���"�U�dAlc{�ѠUjq,��2�"v�����n��>��9���J�C S�V*�:��n(�����������=�����nX���~����?� ��R�@��Q��v<��k!MhHAA1g�����AYS��?Ť
(���*�ۍh������k������B�*��I����mk����-&d %�(ئW6��M����0��\DO�O�yi`tS��3���9�_�ʱ�[>&ΰ�J�Ph$Mw}��j��|����c�;���lC�}W���q�|Jf:e��!�����ꘉ)t�"h#�u������,��bya�&w���
�hR���r_�0_��	]���P����r�$���j��:uk��|g�����-�6����U�r[��K�A�b=�����?5�9l!����0�Ȟ��Q+�ND��Wh�4%�f��"��v��	�o �"�fEK����R�H��Ek�~'��7�q�A�lEx��v�Q�NX�R?cѿ(�0$֘�?l�'�Tv]G��:�y%�����M��	;x���AB���4�x?��n�|k�/�
��.��*�N}�Uȹ�@1���lFMȐ�˸ʕ9THӠCB�L�p{O4Q��]\���˞ �\�"�&� ��q��r2e���hL:0�_Br��X�~�s����Q��pe����g:��
x�ð�]�a��Ʉ�6t �h�ym�J�m���\-�	���Q�5*�#����
�SޗT���M��K�<B	'��kn'�@��0+�b��.ٚk�/w �K�Lr��g1��B�ľ�{�"�od[f�N"`g��{܅Ԏ߄��2fV��ά;IG��PY.���
	^W!�nc�&o�l~�\D�1����ÛN��b�%�ߢ��1� p�WgJ��;���&��h��n ,6���;R�_�k>s���h�L/[_�)�q���́�D����T����\+}����%ǽ�q�����](	"��vh8��#0�y�����i�(v��j�e�o�f�C���PXԾ���b0�Ds�Cn�+6�wV^>O���S��ȶ��V�����է��Ae�'�$�:&�|���[���4_�ݭ�ŝ}/��������9�3ĎA >1ʓ*�쫤�qbR��:�Q[�Ut��j�G�#���w��V� ��H�K� �7z�"�{��ז��%[���UG�f%�k�}�4U@Xz#!�H{��/zvo���v9	�R�L�'��d��
^L���Q�$�ױc��`���G��@�)�'P�w�z�LjLw}JеjM;2T����Iڐ	�Ӭ�U;uyz<������)�����$m�e�ls;�c��ƣ6����1��Y5/�@r�^?�c�x�'ʷyµIW��[ԸD�^���O[�/���%S��a�O������:���p�_L�t�,�%8`���2m4Xor!WN�$alv~�e�~�PLJ��D�t8�c�OP��^��@[���*���U��i�q�̢��������L6��>��Lt��97�G��z�^7�'1�k?�0Z�tT�F���}�+>8wf,2���Z*���:})�̀?�J�������A�����Ψ�^^#����F%]|��!T�Դ�U��*z�:�F�CL3v�6�ǮƤV�?b�VW�c��������C'+Sx��A�~�U�B9�(?qM�;�2�<n�&j��ϓ�WYi~2�>>�r2������6
-��ah�Rz�����9È�5&�����Gn�'�<io��b,D�,U�`��,�,�	�|>�[�o|�����I� ������;�@7�0-�d�],uV�6Y�`�B�.*<�x�8x6��.(���"��K�������m�ɝ�v�u@$��33!ҷ���u�׹�z�]�8D�+��笘�'�:����#ɍ��Ɨm��Ve��~���������^)H�f�X���^u��G�F�����>�B�@L��`8�8��;�������w��R���Ѕ#���R�0�u�(��sCE1�OP.��͹.���r9�)^�D��@.�(�1+�Ƕ�C�k`��rд�v�jʹ�e5�t,2���?�O�P���ڼŒe������ytá'�:��#6V�F.S'4P�'�q,X�pfs8���X���B˔ ��k@z9��)㕽oѾ'��.,��ѐ)+s&����4_=yĨ��9�h=ꓜ����!��Բߎ-�zV5����̭AfP��_]	Me��S���r�@�	oÏ����;=c���m�A:	ҙ���Bz�$/�:�vp�/(�����k�1�=��!�r�	����V�Z�G���#M@�c���,g�
@�#��5��/�!^NH���|�^m,{�����L��^r8�z�|����;�9���v ��>/��'vjʉH��o�NT��j60���*�S�e�Qn��\�NŐ�Tr�G��>u�G/I�<#��阵0(l)M�,�F�L�0[�s}p���7�l��;1�g~g�o�����Q����(��wgM��
�cm�̲�t���a�-���U%|f.2�/|����ŌJ��5�!;���Gcԗ٭
X���A���U4#3��S2k��iK}>6
YZ���9 ������!Jv6�x�	;t�3D�u

X�:sB�ÆG��3^@�*��'��>���$>xto�h������;�YV�w���)�>Z�	� ����TL��U�(�ws+�q�^kZto�#O��妛k���?<q���2_�[�����T���-�� l�Dh\�%�XS,�������ӰGy	u6A+|n�aF�:L�X��2?I5�xZgH ��d1'�vq�:�ͦ8"�j�@� �E�K6�y�m�Tpg�ۇ�q��~)��IeJ=i~�li!�y�w�J6f8�gr 
	#��`]]��Z	ď�����}sS�E� O����[lcҍ��X=�>iU"�\ٵa��y:-P��}^��j͇'҂>���\��6"�@�\hX���n.(���oV�.�_`����@����ك.����Ɓ�4T����݋�^��{/�>���reaI��˖��rb����Gu�jgl��/hO\�!�J����66g��|K&���&�L�a�bH�Ep��$� f�ˆ�65�b��5U���I��t�ܸE1�u��/�+1+�R$h|ke3]��(�;"h�?Rз9���!|y��a��D��u3����S���B(���&����̙0E��c���K#���q�vĚ��s�;�炢&a�}9[[E:.����
��m����*9ު["��<�="�}&�3�6N����0��f��F�O�@��ӷ�dX��#�9o9���ܭf��l"�ŦC�}�#�[��uu.��a����ĳo����}X%c�P_g��+��ٲڣ�!>g_F5��S�JsH���')X���Ңi�e��ҋ���_V3|�������YFe<��ϊ���Ǧ�,c@i�Z#|��fbO��VJ�AU���^�3A�V\;�� �ةA52��35���æ�;/߆���||g&�+n�L���yq����>�����6-Z'7Hbp@+�HC[�U>�>�%va3�P,��;XY3�|e�'>EBf����)jO���O�O�&�SF��p�we`p�eg���DXv3ު�34�+���z�>����z�g���r�d�k���F�a��T�DF�������R��t�IS��~�t8���D�)��g$~�����~�n(� 6Ύ $���s@�4�-��ā�*��u�ۊ�/�d���j��.��K�!TV���L	.J��:^K�JL�{*_y��Ȥ����[M�ܻ75QU����p��\����q�um`� ��*q��N����%#��c����t�{!�Mp�}�#-cd/'�B_�G"����]���O�v�@I^���Fb���x(
�eY�7%X0�{m�!���K�σl�^�k��X��:q`��-��<��ߥ\�|<��w��oĖ�*OL�T�#6���	�8����w�Z2�/B�\����1�o>��bK���������@�����]��m�ֺ(�Da��Z	Ҧc��;f!����c�L�3�����,D$��ڀbÖ_t\���7SD �;�%�������ʣ7W�{��#E��O�)B�҉��Fg��"�؊���Y��`p�RK�?��J�2�(0���*�!Z�]k