��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�KW�UHս�K�7b�^��<{�+LP���E�[��,LUU7��o�9Gj]>�U7��w��L�s3~/�E�����Z���1�"�pK���;L�P�����^��c�f��5�-���j�x:�Ӝ�,o������zi��jWvs����hT�)h�����Ƭ2��|�l���XW��PV�cJB���"�1�)��F4�P��,9��r_�o���!,�!������ʼN�BӸ~���;$��,=��[�u����s�U08��
dѕ��6������Z��gLU�ˎU��ϧwO���DM/�.��j�X�;W�Y]H� ��9ߪ��c�X�Su�K�����C�UJ�?̃��XE�+�}��	���[���C�V��z��!VXNF*�.@uL��Ms �$���t����^�xG�Тhţ�����+x�p=���I(y�D�#���o/��I\����fGuO��Ũ��fA\!0m�Ģc��&d��VN��3����A&���e�m+}N5�+�ut0'�`�$���_��������k�U3�헳�M��䞵�ң�:� �l	6a=���)�`�2�~���]�tݙ���,���;�2f�r>�&�AJŨ!���B��&xL�:��"��F����˹އ�{{�l�k'K��б�z�D�
���}W����K�Z�f'��S��t�墫'/k+p���x&<&�<H$^t��1�蓶����?Èq�8N�XlzG$���W�1&�d�V^
�f����n䴉|��vtg���E�kʦ�لQ3{طY�?u�B|���#�*�ռ�#�4|?������8ccC��������ruX\�LtO���L����,�<���,Zڀ�zh�A4����TD�Z�^���Q�g�Q|�e��3f�.�|5�I�{ݰ���9���t��wA��b�$u��%4RVI.���?�D
��'E�%��������6kI�-�+�e�v	��B���+�KF:-Rȓܘ�ݦi�|,�&�
d@�|�<�1kaJe�-��'A����Ҫk#iFnq'O��[����z�%��{�`�<8���RL�*���eQ"I8�����
r09d2Ū2��XFm�=�����R&
�JI.����DTp�Cb��5E%���q4�}`W�4>q	�/T��E�0�Ν-�P��8��ᛀ����>�#����/Vi"<��"�;�ab�M����A��ն��e��\NV�F����Iz]��YVe?�'��z�E����jS���}�\yk�=1���Xۡ8�P&��9&�Y�ƺ���G�)��h8��2�Ώ���j��WQ�B��)Q�� �$���(���&M���߼B�7�!�n���E��]��P���n7�2�m���c�NԄ��	b�Bt�%�����<�0������X�����D%�������*g�Dn/�b7~Yӄ+�X#)��$�����Cg�|s�.��L�_=U^<q��w�����(�|#}��I¢��t�d�d���bG;�|UQ)�G~������*m�!�={굫=2:�)�B�c&d��LJ� �48&��b[ �uDI�� ��C�;m�<�R��a��4��X�	@�)�S��V�mOi=���'�?���|�0n�u�Oዅ��'�iw���Xҥ���"�<Q���sxN�a��J�}Cb���&FW���p`�N����� `C�넆O�2V/�2ߏѿ��n꽮��������M�ba�}ǽk�a�����~�z<�����@g��o���n��8����~VG3q-j��:����gN� X���>�1����#������{-�f*�)m��|������hֹ���7$C��u�N��f��W�ԡ�Xl���:�'��x��.����u����AߋJ�(9��5d�+����x� �
�c��V�T�8#�c��Ě��O�U~�1/u�Q������d��9ؓ��|ǭ�1�Q�K|��b������6㸐�7R��:���ڠQB��Uژ��kz��,�.ن^*�]LL��x�6����EF���F�U�!H8���_�����D�
b�.}��]o�mp��:��q��Vj��� 4��Yy��g����i��h!�T·o���m]�7����'��T;�!*`�i�	��ai�d���2�bv���Q�� �U��|g��������H�QQ��;"ߓ��sV�4@MN�yQC�x>���z�+� ��h�X��þ�*��N���4<N��&���T]�Cw����T^_��a �i�C�� H��+&;��q:Ǒ@��L*�ﶞfw�6~ΠD^�&=i��å��yt������mgZ����3Nk�!�)3I��"�&%�@ӎz�ðt�[�]JGȹQ_ЇW�3�%8���ґ��Z�Z?g�4�-~��u�igY��X� |DR��S��M�M�@�Ǒ��$"���ch�)[���9]��õ��L�]��*ʍ����
�� ���Žq��6�����){׃~�c#}��$���a����l,��t��4O���"�_.��<���Lê)a�)���v����i`=���e�2t�|"�q,z�~��������4/�C��SR|���Vg���u�T:�uݧ4�6�����i,�72f�i�XV���!G�����h��{TB����~'�R�٘��~�;+������6�����^�s���#�8�P(I�e9��i��N��(ַa�:!�C�A�4haЍ.t�1E����\��N&�1�����6��Ԓ�h��W�'0�^0��вP[��s����}-l (ҕfp�`piWGJxN��!����󕸜#o�	�˔��QaM���l�6�e�sIf^��� �rZ�׸������E`��i$=,��:�"�@����ܛ]���LD�U\cK��v4��OΌr�l�o�r���@z�%��N`X���40�WS<�m�a ����6���xK��O��6�Mf������7X�.;�q8i嫳h��b(5.�'MJ�U��S21WJ�L��f�ȕ92�����\3Szaw�k�_��[>2�q�&���c�zB�n~��Ёދ �5��-�6(�-��0����+$r���q�+���B̝��=oə�qG4�>h�����)ڧn��edw��l������xO3�&���Ĥ �E��r�/d�,��$o{��/w��t��H�tT�P�������|ݲ��ʬ-w8e19�ܴg����:q�HItc��������cJO�:�.��-����=����y>u?�wK�M
�K�E�s7�FEǀnO�z؄�5�I��D O�X�j������>�)��L;Pks�.O����9���[�ʻ���UH��|�qu3�y��E��[*�4�[t��������QGT2;&<f���Ca{&��+' .\4o눦Y�IE�>1���/K�#d�;��X�#�D�F(d�0mh5T;2iF�!@]xZ �/5<Y�=P�is�0_�.^S���Mi�q�
�L�P%�A�rŪ�S��_͑�}�5�;3f�ǩ[�Ҫ��Qx�J��B6�r��7��$�E#N솙$�K�
�J��Y�~����:u��8tۺ��;`_q�z�%{�\��_�뫼�!�+��-�Zp����m�@+��,�$�F-皴�#4G*�u��Nr^xG�[g9��ӌi��ڿ��:�1���l�E�=zpm����hMR~!��`wR�2>#�������κ570�Y}�=f߇1�I��;t�nV9�
����ۦ�9p�w7ڥ�$ӣC�R��y+ߤ˅��Gagc%�S#��/L*�BҲ�U��@�"]�@p�i��EO�������I�ΞF��T�ْ���2�f٥!���&6�a-�Ok ��TɂZj�y7Y�fţF_GKc�:�O���}�裮	㠴��ـ|N#.�b�y�`�av�lX��wkG<���ثc�O��&�Q�eR|Qk{<+����u0wk�M��zr�WC%����C\Y��Fu�XJ&6s���rHm>�2�u'X�'�i�M�&ʅ�����,�C�AN�u���yz���(������.�cx��Ö��OО$���{'.�@����d5�6�BU��-2s\��R�ͣ�j�(�O�d�'����Ğ[/3O*J��9�bi�j���㤸�ϕ��<����:��	`�)e�*�y�"�X?���i}��@�6�����H�����!�2"&`�	���Tg�����z{����Z�W���9i�� �j�Q;�Rr~�/;�}�_T�=��Z�ԇ^�Cj�)}o�����P<{t��I��m�}��Oa?@�2�u H����ZM�~j��\����$�2}�O*����)Ќ�i���/e.���QhMȠ:f:��>s3Vpþ��o���eC��OI7��6��#n�M�"��6G�r�&�������$ھuJ�L� ��S7,	�Nt�L��wC:������{����՛��g?G� �L�(��
���ٖ�VOF?@�@�>ɣ��)��W�T7�r���l	 `hw�y���J���1�OG<3�j�@�A���y��2�+��$y2�A>&�O&�S�% ��L#�VÑ��Х��o�ֿ����4"c�1ތY����>�T�~Ԉ��'�G[�U�
@<A���Q�}�j +��!SW*O�g!��`h}���x�ٞZ	�=՚j=��H9�6�zD�:��j7�<p�;(+�����S�6���=���<�6�P����(�ivS�4.a�}��O��N.Dn�^��Wt]R�1�%���Ȧ��b	��p���Z�'����q����A�B俔'��T�����B�!㘥��A����)wsGE����"^�,e�5A$`����a�e��`��K��������QV�[�gW\�E)�Ą)�p�i�Sky'�j70�\����VM��c7��LqD~5=pr�Q�gA<�?q�4�i��M�T뇫�������	�1�kq&5}F�����C�u�m�W[�m3j+�8��êj7�>���%��~��-/n�)�������?�W�/�Z�/��xм���H���w��M�e����.S)? �Y���簾@6H�����衐��Ԇ����q�[�n�b���8g�n��\Y��h�WC��x�FND�Y���:p[S�C�t��Op7%H���˙�� LH��S�N�#�q?�&����-jm
Uo[
(�~�w�BxRĄ����2r�-��l��?X�hm�q6�~R#F-�g	�zR�k�W���%�ʗ�j����㉗2�yGg�8ެ~��a�r줞m�����y=���+�_m���ګ�\~[vǊűؓɧÀ7�7��*W2.�wq�8��=>�ޖX���s��l8�\���VT��]B�m�>��c/XL_��a%�̗���,�yeه��6$H�w�NB˵�p�.�
/ܢ��ވ���M���>V�M����Р'P�"�JXS���J�Ͽ��+�Ql��)�l�]E5�^��.:��0��E�c�'h*�������~����ZLu@�89b/�_m%�w��C��O�)�qd	��Kh�mjBEh�]
E��U�Pb�+�zȒ�죤ۚك[
iAP3o�$}P�S���Ԇ��lx�dd�az����~���؀J]��Y�ɺ����"��ڷI��?{�ѷk�8���{':�ռU�z,Fͭ�!:� �l�!�Pȡ�ݖ]Uy��\�E���aN��2�����(B��P(l�	JY�;x�]�7��7Fo�>p�$���lc1��� �F%�Y9�5yu�1�w-Y%ޫ�"��T�6vW�(�el���,� _T����ݕy.��U� �l��]��	�@@��o!�.��E@R^e�p�b���!��@�PGs'��
�_�X���nԏ�slz�16�{���=k��dL�������8Z���N
��;�4[� "e�Š���!x���Ǧ�����DR!�U�3`�3⨵��n�[�(Q^����5��(.�OȆ�l=�iF�?���R�̪�;PB�7$�{u��Y.KU�wPѿ� �����0��z��A�[P�>�&��ۄ8�Kl�(8�=�S�����*µ+
<�|�Ș�L#T�7�֟�f�fü�qF�1��92o-uv�cQ�\�X�c߇��C�
nδ���y���� ��#^"a��܎Y��^��H��c�?x����-�J��4��:���>�6���N�Y�8�m�1�y ���'l[w�w-�ʞ[���Xi���ϫ}*0ckR�C}����R�;=��iq��X^$�0+�wBN�����T�dIȂƫ�cV�o:��I���W��L����NT-�F�j�?����_B$J>#Wr? � �C❭[c�!�ڪP:�q���d0��xf*��9�CƄ�����Q��T�aM�7���|��F�k�D.�4��YXEtw�����껵CY�_y��y�|�zPo�F1��SY
9P�x�������0r���9E(�U���;�Yb�K�T/�'��MP�7'�)�L���d�Z�f,�F1��4��`�~q³Zk��������T�0��=9�i?�y�k�q�7Ĝ,�0�۫�� �K&�4�18���6�g�&~�J�9�	/2���h�Y� ��Z��(��0�j0Dд�j��ڄ���F,� _�K��	⛽�4:&?��.������j	�k�xi!o��h�h"�*&����{u�9��b�� ���試�0�%���a��;�5��?cҤ��m�1�0�#1+��)��o�*�v�ߔ��m��ѱ|J���!���Y�
�X2�n�S!F���]�Gu�5ھR��Ң_z�:��K_TBH�ȱ���w��a�3������l��ᰣHV\���'�����Wc6tۃ�>9��O�	�]��C`�Дq pȵ�z�'p�U�����t8_&��n �<�k�J�g�h��֒��[e}C�Z
;��ǣ�t����0��A�&� ����X�'J�WC��Ys���f�;�ab���l�K���A-�@[��U����WJW�ɶ�O/ǔږ��H��pm���p^K5�����x��t^��Z{��8Ql���Xg�.�bt������2E��6=X�4cĈǋ{?`Ul:�¤�D��|��+��uP���x�5Ú��8M��`p�{o�K���Ň��������\X�^+�'zl+k��о��B��V�h��X�%��tk���N��@U�����)Gy�d���DW���e��~W����˃*��]��b;d)r@-΀�_�q��W����*�A�o�TX�$� ��%P�$�E�r{��C�g��=D�59�Fí"�^R^wl_����5M<1t�"ak�z������o�	,��	�H�rElX^�4�-�>��YW�;�5���C�eKNl�N� ٬��wWK�.D�R�{��B!]��dJ�ڂ?̊;(��o6E.c�B�r�!��?`�|���'�{>tw�@��3wO:�@n��CPmBo�e�R��°V+)��#�l�}�:�{����u+�#T��klW�7�K#F�h )K����,%�Of�f�
d�ZZ\�j%��$�yZ�RW/�+{|I���X$��ƭY��1���~ū��SjT�&5�+�H��9^�����be��YpQH��+�>�^8��"������(5����x��?��v�m�`]#k6,�/�!���.]pt�f8�hԺ��{�J |�ݡP�������`��ᓴq��q�=��Tw�a�6mɼ�E!jLd��߈�N$�$���_T�$EL��4�uuN�PIIO���k)� �����c�T��	���1�w�Z4�@�c��X���kZ��>�5׾�@�g�����'-�Ȥ���9(������i�k����u�-�}WĦ���F$��~�6����)x�{�4���7>I�k�]�>	KZ��x�OD����� �<S������=ڧ�2��E�y�-d�&�/"��Rh��ĴRV�����2\'�ݭiY�!��Lk��b���#M�����B�����J�4���7�����M���-�-B����ܭY:��ߘ����ȿ�8�;���6�%�@MT����C��jZ��\Q}�6���Xo7���^���<�.�>,�}��������x ���$���(�y�,�&�DH
�"��Ŀ؊j+u�G�#rM�g�1����tZو�g݁뗖�K�	���8��=(�ڐ��I��������>�8�^�|@�դ3���N^(� �%��u�ٱ�I:��4�RN= �UVb{��� �sD;�p2�,d�ae�m�/i��1>������9��{�ڈ��b�Un*]C���yC���ھ,:���CZ}��C�z �v���O�~�ƭ[����L��mq�Ծ\%����ϊ0��*�8���G����",��*ۜ����x��g���e��Q�a]�7OVN*�.�a��uh��y*ځ�ܚ��D
6ګ�2&m��K�
��a��y���A�K���"t�!��Q��"�W��
��l	ͥ���W��gI��w�:��0:u�I�:��漇��q78�T�Z�}����v]��ܽ��{�A�'��fE�' �JKq���Ŵ�t�ȍh÷��N#DTb�X�.rZq�ܥ�p��-"���ɋ���}� <����~�Vb��ǷR�2 Oa8l`�F�Ռv[���e��:��ң�������۵����3��N#nKo��i��%�[1�nJ�Sc��.�-��#4[ �����S�ҼA>J��E{��q	d����$PCY�vqo�L�ky�d�=B݅�9q*[�:���O_	���}�`��iD�7��}hK.���rp7�BP�k4�:Y�ĉ��մ�Z�Fj�t��!���3�j�P�Z���_Z�ht���L�!�j���~��)�[C�.)V11-Z���i�����^�֝�9����ٮ�,1�\�Rr���Ԧ�
���i�ɛV-v��(��5o�+,Xن��@�D�]���Y��y>
�~r�3i���Lݘb
��¤��`er�_��Ƒ�s�1
z�p�٣?��$���cjOü$"����/�׫I�A_��T
 ޴�U���;O���	e�i]�C{�
?��T�}������"�����c�G�K}14���i��@N�_�5���g�h%.ԕ�9eٗ�l�^��iW������|$�&i?6�S\+����L^nVh����Wޗ_�"�k�����޳�ET4x݌��%
L~��d�*܅ ��F|w�`y�j��e�W��t�����T�⌍��D�s�?Fv�q��jܜ�V�������Q0����1U��
����&�?�);������W%���+�㵹�*� E��%�OAj�x�+�2��|	�D�plO:�wS�����q�1��7Nu�������=0�lb�?���n�L�M�w�;���=~����+�#~?o<�ͼ��h�E'��*ۀ=3c�6We���i@�&�!u0��@l�R0�ָ����H�I�\@;q���6Ι���J��q�9���<V֧��X(�Ρ-WF`��U�����aw�z<��=��5�@*�z!��8z�Į({N��"�Η���&ܿ�NDQ�m����&,�b�� ���8��Sc~�|w|ca�0`��n�2O5o	��o��&X�-���Ur���	����MD�>�SZέ6d3���St],����!֖
����7���sQ�^��%���Kg�a��
,H���[�W�a�:Ђ�ѧ�g��.1Q�ϓ8GF$I��g���;���X�l7gYe��\S���K�]�ɬc���M��	�,�4��U��7H�I��Y�kP�ORr�$gs=��x}��b�)�N��iA������ ����
�a���PD��s���4d�*Cˁ�������4���s�j����bmR$hva��<�Wꇉ�y�mZ��\�#Р�n��k����$E��|�V������.��.���t�\e%��3ي`Px����r<"�x����O�ly9�+��0��O*��+��ZG���b����}�W8.~�c