��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��ᕫ��H��gq�f}���+����c��0�7�*�y�HXH�+��Y�Ar�#�<�k���bu�-��.���O�;����b���7pE+�������v@��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾��"o�x(�m\񗟅�:��e��Ӌ�~�fT��K����O���<vբ��`\��t�;��v�%&
Y�=�2�|�mY�"x�VƱ-� 1x5�f-�!ԋ���K�'��N���/I��yL����w�뮦fGLW"�"���<���1 z�UM��2�H���T�������\|e�B�2+�����i{�ΨS^��'DoD�L�p:��@F�
��2��ee��i'Ӹ#� cgem`�[ ��P��B�L
d*f���(��@lS*9�~,do��-R\rz7W����� diN:��l��p�!`�qN�G럫��Srժq~�mye���q}���5UI�v��γS�S��^أ���1��I`F����>F�ϊ�Ee8�C���Je�:5��r�ż��W_9��i7:R��T׿�6� ��f�4�`���w�p=��⨔�J}v�Rf�*oD&�?��K��,=����7��C�T#�5���q�W	�-�I�/9)af���:)�������)��?��X�5�AC���S4���\F��;����o&��%�y����J��k���!�%�wS�(��?<N����FB+�q��jB+;�� ���=��Abdy�v�Y��R��9�|�������_�/�>N���H�,���+7s*m�,��<6�ǥ��� C�O��G�OS��`�@���$�J솨����kN�%��Q�r.�8���2}�ڛ��mi��/ì����|H��y�>F`s�s���o���� �u'J�'���N�z-��@�x�^� m�s'1f=�����/.�����YoEp�=��u�ɴ?^��
-�أ���h�,�����&RWJ��$��K�Lk���`x�<�vfo|�/{��[nʢ�5t�����/������I܌�Ko�Y7��=Pʞ�ݲ�^b+����T�4��Xɬ�^&d��b���?j�80u��4��&:��J���޺8]I��ɤ�"����w�,�$v����(t��۬��9I��~�=�mԍ�m��%K\v���_�[��x�y��xm��?H�.AN��x�۔L�S�2�,�&d|K(3��aN�l�#��cg�����E~�>�!5v��~���{zv_���/M��s.J���AH�О�K׉��T�N�bT��\��tv�2�I݀��.�Lt��xV:twÕ�j�v�&2QA�DOMB�y�Q�꿞�- �n	��������85��	��Ϸz�����ƣ2��p|����&���z��X�FS~(&s�Ƹ%.i�æ�F59$�"�#�h�љ��z	���,,Kɺ4������k�35���ј�q+�JY�a�HYX��F{�J>�s�����xK���	�G��r�D!���U܏��Y���!J"g�:�}����ى�+�ؚ��C�����,J�����+�xZ�x�����nY#F/��j�j7S��U/Υ�}	��b��~�PT$���Nt����7(��1X�a1�!����6F<�E���ޟ1e�0�|G�S]�V��k��8�卒"�o|]�������/������o���C�%��"��1�wD
���m\�@�s���� ~��A��ɹۡAC�׶@���R
��hm�
�� d�A�IE5ע-;%����j��r �Hfw9k�E7.�1�~,\�v�USq��ޢ�8sݹ�O>gǬ��w�-G��P��ZR-w��d���J��r��&}��e���e>)O3���5�>����;g�ʹ�~4l��8�L�~$��*@�̣ޗ"��3�ʠݻ#� �OF[\F��n�����z#�Ԩ���!�,4V��t��y E��P�����k�>�h��@3�;j����F��}@8r�&.�a�^9n�]&5�K�Ѱ4�5��,[��0�-63�S��ϟ��`���i�WA�����SN�|��I
��s	����ҽ��tFB��VT�5)��
�<(���C�-F-&��(p��S�R�[%�/��=nwM�S�F�H���1��ѧē2�J�2�!�R�cj�2h;�f�9��5��P뢖 af�a�C��Mt��	Sx�Z!S���敩���� �0�̣+qs�p�z�ߡ�z�N@�bT:^��)?<�./Y2�6ٿSb�B�r��w�C���ϏO�b�ܝ2&8�ȁX1,Z����dA���>��́��1�oCC�'���{�M�Wk}�V���u�FL7_u�A!� oa�=��Ռ�F��!m!d_�Lk��2�:߱20��D���xX�����݃l���;�Z;����"_��rC��etN�l�%<��q(�Qa���K����7"��Wj���}���s�z�ײ����X)� %S2G��@0;%i�V�C�F����-j���*&���H�y��\������!x��$��kn Y�J��;�֎�>�'�@
�=r�]�Y���]�'(T�wLќ���λ�p�щd��H�F��AdSl���|1�cV{�bd� IԳ�;d����Q�ݥ�-\W�>�,2
bqQ
v���K�X�=?qT~���Ջ����N/�b7C,�/c"�=FԄT
QF��ݣ�N��.%~k�F�H���iڇm_��S��]��2�R��C�+%|	�@.uKE/��fŰ%�X�A��(	\�Ǚ�&�K?�_�7V�3S��gc�n�V�z	XӯK��
I�3�Ǭk,�&�������j;�z`�g�\��"p�Yڡ2��Nz�};��t��x,PYj谡�&�J�M�wj{%1E=�x������0 ?A���e�6���S��V�T��y�w�+�F��`�&��l�ݹϤg�]A�`(���>�V��VS�`���cf�a@�l,L��';c�x��P"�h�~�����#�l��>�z�Z]���㬚�@i�c�;�}�%��:�6�T.t�7��h�Uj��V�&�j'Ϡ���CQ�#ּ�;�fq�*�>{�������I��~�q��9�A=\�������$�h`G���n�=���q��i�1�ӥ|XDG�J����q�y�L*d+�o�������v"?	�UR}�9��3�0(1>!�H{�B���V��a��hz�ٸ1]�.��1��Ɖ�\���yid�r}�{�S�UIL\8�G½g��ZdBTQ(�g�M�@(���=���*@�[;���S
Qbd
I�����[�q4_)����꣭�y-�U%��O��Z |�L]2Xݚ����>B�-����g�@}�Vw(�#�J
s]�:<aˎ��_KT@җ�o�i��h��PR3AdB�;Zѭ��b�h Q7�1��S$^[Y�/�f�gV1�ŌC�Q/zZ��.P�L�O0A���RX<�tF�f�`�m(2|���!�����?��Y5H�>��������`s�T0��X��`���;h���<�[au�ΐ�-�=H�,�P�q��$�M�o뀒�������}Y�g�ц@��*%B9	}WΟf�E�p��:��~g���;��(��l�]�M�׷*���e ��,x����i�K{��r� ��D�Z���wUoR--�[�Z@�~����)P��ُ
sϒ��nE��[3�ۂ]���t���7&+��-T�"���0����kQ������noA���e�t|o��	���t�rMhG���}��I�����ضNӏ�6�ν �΁WKCL�[�<XH�=D��|t9��jT���ı\��-{oR�Q��)�ׅ�x�"NfNY�e�6��(?�~�L��_��T(��p��������C���K�!�6/O��v��Z Y�3���u>%Ͻ�9��G��E�k�'u��9J�uK��c�=��&V��p��� ^��4ڵ]Yx]�u����+u�FG5xw����U.�)��;8fµ�l�������wr�^($q�� �F�	�����}�sؔ�����,����ћ��a������UO�>��?vȝ�rW'+��q��D+��^-x�>��Q�v�$�
Lx?"&$��_�ڀ�b�?|)���琌��W�P����y�N�Q�n,�z�rg8Ě�@/����V�#X��f��v��t��F%q�obvYM��܎%��н�	�M����{k�r�t���rEP�>���5�[_#���C���;=���z��i����?�Lo2�w����*k ؁�:3�=�=��8`�`��Z��'��5���_�����q��OM��Nc,�:%Q�$jp?T"�p>eL���b�g�P��_+�3����@|Ϭ[{<�^�!%�"�5�#5������q��o��t6�' ��i��&Z"�l]*2�8O�1{7�s|��"68�v�����c��s����H�Hl.{T�s�~��]�)�>�OV�ji �d7e���?03�:]�q;�\Đ�G't&/ ��>r.<	b� @o�@C��]���6ha��X��;���2����
��y��)^k$��l�-Xp�ו� v�}l���į��ie�د7��'ɰҟ�C��|�^�BrSw�}˧�o��u�F`������-�ȣ�V22�RF�?�7�?�����3bHy-�z�����?;���K�j�K��vlE�^5`��!�=����HtSI=�x��_��]�%P�+�����M������1��YHc��$^�@��s�|�l�p �q�r��~����3�61��%#�a���m纫�4�D�v�Pcm:@$���o����g(�����Al;�N�t��A �Ra��#C{*�]�R,UMna��1F�(H�f���zgJ�n-��T&owD����W��]��
����<�+��"����j3GEetr��䔽�r�
k :��4ӕ�i�f��
��U]��������*���50/�m7��P[����?ڔ. �2�ԳR��oҡ����E�Nh�Ej6_�Jw����f/�ۄ�e�=?�^�&�-�8f聞�o���I)$�j��SO�(�u
�6�$�v��C�á@�h�."�9az��Q=u�w��3�d�}���	�֜s�� ��@=dq�.D�l����O~�W�X���6vDR�vz1hf�=_�Y+�e��^o�9v�篎a!ݬN����[/u�C�V���o�5��U˦r֌���ٛ΅R?N'��5 �Bz�V)��������Q�|���aߔ��x�*�HY�stV���f:]�l�n�e��=�Dj�Ad"Q(x/�?��U����۴(^��=5u$%�� [V$�����P�Z}j>�{E�O�Bel��x�lU��/�A%<���y R_��}�ƥ&���}
bN�s S�]-k	�h���h�>�:B����ы������a��n�g �����k���a��"̷��`v�Lczs�iM&{ 8;uf�8�6�:����G����R�#�~�[yӮ�+���w]���X:S��g�ܖ�f}0�P2 ��e2o���8H��Oi��M��c&�Q��&�)k�%(W�y.�S�+�Z�Y��J�A�ז�!�X#B5�������M�6�"1p�A<j�^�c�p^��1ݘw�j	���j�j|X�'�ȟ`�S���4N��B��pZ�}�$FϾ�;�~w�ACY�ѵ��6
���7Ѻ���?�uo��Ϭ1�!V�bn.la��ɱ�-���[��ĵ�a���$zR�,����L�y�����L��i���W����5#f��z��[�e�W���
Z��(��͖���
s�%� Q J�/-���=�3�pNg���|��n2Ű|
m/(�d������E���@�<�s��iNywC"���B��V8Ɠ��zT�L�#jZ��ٽ �����?G��*x��Ц��UW5�L
�yӒ��Q|C�́�+�ݕ�<��T.C�'�'��S�ds�U�)��2���U����n�UIf7\v��4�����U?���"��	o�bV"��>�ߖ10��s����uz#}��ꙏ&O�=?�~�D8�Us�)��|d���A������3_�%�W����b޾Ǐ%Y��"�E�![{d��`п�q��k�F!��w�'Gū���'�+3��/c֓(�X!2RQ?*Ю��2�;z�'�օR�� ���ְ�ߪ1V+&��5�uﮩ�h�R�� e�v�*%P��kQZ�6���p���7���͊ķK�=W��j���{&ɨ0�=&y��x�����Zp�R��:}X2bͷe�����6gHQ��Wbfg_�Қ���%ҩ�-�'ɁID����,	&�0k!�oK@Jé���F'�Wm��.q�2fJ�z��%Irl��M)��=uVO�s|�m-�}�N�ݔ�r�
^� �w0ǥ=,��+�s��Ʀ޶�e�B+�;����Q��AD��N�v���ݙT2Rq!���YK|4׀O�bu�Gҙ��RqgMp��K6��x+�"YƠ}Kݽ��?���e̳[#�$M���5��}�mX5ٟ=#y�����W2%mʸ��;Q��,�sj��S���I��y߃
K��7��nKp�$���40��5IR�.]��K����lD��?�#�M�D���><�?s�ri�/O���5�;�1�S����^Y�_37��u�Z�d���n9�49kWj��-����4_�^�e<RT�S � �`Ud���ը�
=��f��ѩ�S�[h�dܨ�� R7��)뱕h�74d�3;�U���`���Ўz�e��~����v�"��d�O�����#� �)QI~� �}AO�I&�9��s#�|��3#�l+hA9C�rپ����Y^�wI�m*��	 v@�Ͻ�rp!�lNͦ*�I(�يdjBB��\��c"��,�-�e���?p�.��y��0�@Nw��mh-��)���
����<��� ��,�21�f���Tt\�����u�2+i��#���"/Z� �im�W���{��~��JO��ZNAat�e�,yK�	�9I�L9�u�1	$�'l���_:q��eQ*�/�W!J���dU|x@s4l@5Ք_@�m�q:���Ww�~�ѿZq��X\2�����{N��:'q��i�p��G3�n��c$��+ԂHo+S �BrY����ҩP�Qy���:D�N}	�k��ћi����y7��$�4�S:��2�2wr1�v��u���s��-��a��t����.R�V�XD���$T<N<B��LW�0>��ԉ�Ƃ�u&
o؏\���91v�����������9�g����[��+�X�QȂQ��.�_��!�}i��O�U�i*w���Klқ_3@�����j"k'���q5�@-�տfl��79+?�ڕ2:*l��rC�z�sIB�"���'�ּ��.�B{��������UA4Z�ҭ��=��щyYUE�8��_[�)�*lb�W����hfnS��%M��Z��?�>�����mh^�8�R(c�˒�:�zq�rO (WM�y���(�xP���RU�Uh����"�-h r��ì5&q ��!m"H-���RZW��&tn��8:0���%��T�s\�}7���g�|�C����t���w]�pa����vy(C���7'aRϊγW"�����? �?V�p�`~���k�i�a���d�&	����Ћ.�&Ҽ�/�ZO�����ٗ��=O���M�N�h�әj<0���	[��r������)Kc�-�R٪��3?	���|��r�`<�`�D�K��Q�uХ��f-�9�hs!��r#]EI�8#�G����-w�J5k�����(����/���j�r������R���o�8#w�7�VX��'"����)L�k"$��29An��bv���Ǭ�%��z�\����8��1T��3��@��1�GS�����:<ɵ��<�k���Q9љ�/'���%o��������Y�P�A7�;Z3���~ܛ�)��ی��7�}m�c�%5�G#���2��F���KP��N'�A5S^t�!H�
T��L������Փ��P4�/MJ�s�[Ы�fʡM
�&�6�m�|�R:62���IY��{�MWu?CE}O�gK�?jBta�I�6,�2N��t�A��+���'�=�����ZjŹd)v��}��&t:����Hn�������%�9E_��(�ڏ@H�]"�$}G��9��؝A8�4�:���u�Mܴ�j�l�z�:�.kęf[�"�:^�J���1W𪣫a���י;�������$3�d�,�	�oq�����
s��x
R�
+��X#uA��_;���Ɔj�m�����``8��c��LoV�#���!Cu�Kיl(o����y@��z�@}0hϳ=�7�U$Y��$����z��2�O��ɢy�"0��==m�MItQX["�� Gn33 L?L:�>��K7�M���O�&�ϼP/�~4)��,�lȔ���w�y�f^����f�c��;�vЬ:�{�u�G��O@���3���[�Z���Wu�����_��9�U�
�[p:��]�����%�GJ��\}��*\a�4��m#Z�#.ʀ<�v�]u3ֹ�ۺ�V&vg�3�!�SPX	������,�A�E6��
b0�R�1ƻqT ı4�qُ�:	���ܙ(j������C�)~6�����@K�v�ܫ�&'fw���Q#���g�ɉ\�wH��b�������x�g�p�}8���*_���[(UN��:ӹ1���2�N>���"`2u��P"�V-b`�)u�X�ċg���U�3Y�����U�mո�3��bj 6`���60ĹX����4��G�s�=T<��'���ܵ�%4E��̓Pn�F��Jq��K�W�Àm$ց��Z&��[ ��ˀ�T{t���!����;&.����Fs����ai|na���	ϥ���]�<R�Ù�k��c$�D՜�*0��\��0�t�8��m��W�����Z��e�ؗU�'x5K-�0�xt�7v{�<2���Ԧ�Q�):�Ds��p1<��L6D����Ml�vɫ�<���l�d��s+kK�j�l+5Wa{H���8���U����m�Y�ٍsnGi��<��ڎy����V�L��V1����*d��(ޑ�)������0�s�����G��w�Ԝoaq	m�t��ZI;����|�6WxAӽ��W���c�?d/����CKd��W�k�&�p|� >�E���~�yiʟi��5��"�̃+
;��J�]R�[l�q/�P�LQ�+���"�r�_�c߹�	;��KE���k� :+y٘j`��c�������}EoM��-�-J7C��o��.��ˋ�K�Fl�kB��{���9;8���/�ev��:�\紥ec�e����'z�����`���w|
�&Cv��\S~���S:�,z�X�$�3�gI����^{F9g����&NֶL&��\��T-�ƭ��r�B%��,�x��͞Cp�\U"0��>9(��r}J��ݸR��JI��Ni۶��P/�{�y#N���|>�\F��2;`w��0{�,��ю5%�6N)a�@���e<	S��M�X����Wz��'%�?��c#h����x�m-{Op��9ص����;�f��Gz|�_j	�X���m-�T�b����w�_�GV�����Y�̨���r `L�N(���8�4J/��߸���3�>2'c;�
b�7"v��J�t]�ǠM�.���5��-�Ǜ��}r;(�b߯�b\���_;�n�J5$������/ӿtW@�b�-�{� Q��b��=����'9ܕ6�T�.zشs��D�2�=0_qW&��
q 8��˝vw�i�L+^�z-Z���F՞+9�v�`;�ǐOu\鍕�kH���K#�\�w���S#5{�;%U�8���|�j8���MA�X�t�aUH�٣A�-t󾙉����(���<!��)П���h��L�oT�%�d�KF],I&vU�sT�g�6V�>��`1	;43;MH ����G�k0b�&F���Rs|�x"o�`����]%���r��X�][�_B6��
,��@W�Y>+�7S��qH�q��dD��PÍ�]��q�;/l	K��߸��-$����/�kZx�����C�k4�Z�+��ٌe�J*,��"^!k�=������>�}�.����q��5$L=�GZ���'0$����H������&�ۙ��u��d���E� V�/���qWg3��J�#F���;�\���\n� 8�a�h�<���<M�v�B n��L����emT�"g�9bI���6�<�b��*�N*N�Ѳ��'�{J�?m�\�YNefE�?�-�R�C�֊�[��K:�Z3�L��*e_����[�_K8-�	�$�q�lh6@��U�̫v��*��ĽI�	�����۩� _�4�|�5T�qk��0
�4������4������꧐�r��I8�W(�∋sZ�-���,�ؾ$xF��7�E��o�L/e�Q@��vN #,l����#=N|����2�&���F�j� ������[<��L���~˯�-��*�L��т��+9��c�x��(#O�����ԋ������
��t ��Y]m|*yB9����f��J柗?�����č	W+�B0��tf�y�Qೠ����D�#��_�!CHA#=��U���(��X2Y<�-�-�.P����֖$y�������P��l)Js���Lf���e%��l�E�ˍ�D��3��v����X����I�A�k�*?��w��𴖺���I|qӁ�̯�(o�H��&��&�q�M�!^M��a���MD��&�_���'�Si��C��!M|�Jj���kZ���@!��a�ԣ�dcܾ<�;cbW��rdx�Y��z�@�{P���sӷਞUr�EY�J�ۉB�\����9L9=EY��<��WFg	�
Ɂ���D��W��;��;X-d,����=B2�Zc�/��Txk��� ��z&�u�Z���F �&���I64|�e��\��ݝc�T��C2�b��vDv���u'���Xf���efY�6 ���~��L�$���Df�=��Od#����x{��^k6(��嵑
�\�3iҚ-�Ú��N4[ا�T��^8�>qaT�Z}�����R&���0ʠ�U)�
��N0;i%E�4�7Hst��K�L��[yBY�������E���/T_oY-�����y��Lk�?���}��9�
�L���b"͎�Ѫ�..�	��0���Ex���B?X���j��X��b��n�2�}4��u����|	��	Ģ�a�3>�m��8x���$d��V_�F�!���u~gW1�蚪�W���p]k=�F��l�.�����W�� �3��{V�ˢW��+V��%�h�{.�α�v�ʸ� �m��w�3h@��T�#7v���sU�EM�NZ�W�rKw2'��'"	�>�Rac�O1�E\
��9�`qx>����\fYP�cO��Ys󭞁w<\䂉xŷ�'&sU�
��5K��f��F�lY9�y븪s����n�dG�K����3�O}4͕KU�4w�y�j��2;���]�՚~�T��n�&�z�$nRݛ-F!"��R�/��;�U��5�9����)����j���a!�jo���<�/����a �X
�ȟ/[)x|p^	/ )38k���T�< �����5{*�ߛ��A��a���/��K��t�paZ���d����R`�%����i��g]Xa��l�? >`���
�����ѫ&��Y�X�����&��1ϯ�լ�3��l �𯉴���x#��L�=����uT���� ��E����e��JYw�8g�[8��0�5e�*�CLFdb��"�(=#]��&@�DP]��"��@^��ĺBcw?pWC�.k��&1t�A��ɍ�b˼f.1�C�<=�dŢ�jyJ�����,1�Ӗ�J�r:l͉��n=s�m�m��B QM$���b(c����]�x"^�vw�i<���>��\�T��(���"�x|��p�*ݑ?�F�[Ɂ|c��,�?����GPX�V�U6ov���Ϥ�Heb��#�q��I|���:��l�5dH^WT��b�B�8PN��W��Ięs8m��fEI�ۑ�QOY�ދ�C�����٭g����t�b%�t�̸�� ?�⾝e���3>H��=��}�r?��mVE�׫�W,&qca�[��X4�;��A��Lz5/跕���\K?)Iwܰ:��tN�`��ʝ!\.��_�B!m>H��˾K�o}-����~1���0$v����r;P�qս�A�7_�sr��{�w�N�$O7l�[������3��t��F�`���� �]1�p�^GP]�it�������!��h���s{�� 3aQ_%'5~Cd��u�Bp\�ٹ��J �w��{Rcp��HU@��MϨI7����g��^�ʯ�����;���T:-x�)k*�[w�������h�q��c5g��h=���C�(�H�i�#M	lz�^��k.1�HѬ�&�Q"JD��A�R"��pd�*�����d~�]�����S�WC�.p��VV�E��I}G�]ݒ��(�Y���(I�3.Cjk �3=
 
����p�t���rX�F�*_�ͱ�
��9(�
�'+�]� �~���u�no�� �X2�#���~�Z�3p�����"9Ġ%TZD�"?��_~H�?H�+t��
#��q��CI�0�If-|�%)�OnXO���� ļ��?e��R���z!)�nس�W��`.fhI,G
Ķ���M����dvINx�{#�x�U���o�~�tU� � �,*׶F��Э0v�f_�U�3��xMh������F��J(T���:��/Zȴ����֙��`���F�����A��)�P�'��/���z��8��ȳ{��G��ڷ`�HH�y�56Z4�3�V�l� QY���љxd1
�2|�I�%���@�6����ؘXn�����5��>Gl1��k.�_v׳���S�2�%���{L�u+�ƒG'=��b{��Q��� %L�(X�ᅲ�-�'=��׾�̜���(y�<fY;�^Ģ$��@:o	ҋ��<g��D}ZI�T}r?'����	�C�J?t�θA>v5������ P[9�^:ApH�D�E88�G�2����`��uk����dx����E���r�C�rnhL���^�D��i~��Cj��n^�2d�����6o��6 Z���(�zpE�&..j���Ϲ���+�"�����?M�_��|N����`0+�,I��&�_�a,.��i� �Eb�����.���m?/��t��@�R3��3%�s�)C5��Wݖ�l5X�������{��I5̍)u�|����Z�5�6�������� ���n�e^��]?{&q������Ó���W1�^#��'$� ��f��V����+ �e�"d���ù�"7��� �/�L���Gbu}�|�
7���������>�]�dl״�)}���D�-�� Ԯ��pK�w��{I2��bD�Yx�p���W��(��uf{ �V
�L5���Aq:n�㒸ZJhPLCG�@�$��)�� �t�M���uJ�*U�ø�0�3$��\Y(���A�)���4*����#4;�6f$��Q��=*��4���D��XB�F�̚tW#�3�k̐C�`�C�S�D�D��V9s^���b׃�ѱY�w�*�v���k	�r�cc�����{s]X̈b�갤��}�5�\�y��Һ��'~8:���x���q�)G_+h9�~أ�NUCB��Q���eB�ksL������?��w0�:���t�$�x<ƈ:	�`,��5<�*Cƶ�Izo���.�(�,��s�NԺY����I�}����:.��x�v�����H�l�t�PH�IK����� [�TF�L�!��ʎ+��7ʂo����ԃ4α<��r�	q�#b�K٣�B�niɇ��&yF�����}"�`B��gޱT�R5a�Oi@i(%���	M�0F)� c���B�ry��p�2����;��X@|����%�o��H�����T��m�i�قÇu�)��nس9	�.��?�;^���X��Z��:����C9�����N��4��L�r_u��?��X�-�ϤJG3���+�O^�A?�p��)�^ڇ�}�r��+��ScnIf�*6����Z�O�_1t�+i���ra�Ę��k_|���>��3�M��Eu�[�ʌ�@�m��P��zr I�2FY�C�9i0%�{�T��Y9H3z�y����0\�T���,�#+z�mdD�9ͫO,���V���f��/L#"��~�n��#�ch��jH�����8=I3\���%feM��\$���-�:$�P����9*�0g娹z�U3Χz �P��g �lA;9�6y`{/�`�3�LYkZ!��L.��Y"v������6�ɵV��'/����8�{l���f�@?��1�l;Zdt�c���V84�6�T:�L��l2�6Z'�����HX�divaK���አp��Y[_��A���+$/��c[��jȟQ�b��VA��$�T���V��8a��oy�7s��W �_X�L> Y��VHK����=��2��\��/B�����8-����B�FRl9�|j�*A�C���>�t`W���|�_]<�:g��
��I�sLۿy�[�xc��N�Nږ�����ԹE��쑠����Z�ʗ�K{j��T[t	�=�`��d)�wf=Fc�2q��Q8���c�1s1Σ	2��y�Ⱦ�G����xr�k�C$71Ģ]M��~|q�~�2�8^�T���X5�z�w�x��B+3��G����r
���cseS�ۮ1�0�o(�\�Mc<F�r�5mσ����D�I/�w��t�c~�&=��L<�T���y�I�⿁��ѵ��yQ�A#���q&$�Tפ]tV+4���4E0Xm�h�<R��[�Z���\o'ًQ!�?4����9)�JQu�߅I!�h�{�D�J�X�2!V-6,z�D�c�'5�e��(I#qYS7�q�ԩ��a�6�~���0 cD�'t�u�D�!xR������]��S�K+��~��B�rNk5/�9�hMw�u�f�u��K�e��7w�>�-Ԓ$
Lc�C�$P����9}d��˓��Vn����X�[�K�Y)�R�[P:��ڗp��3졀!w�b�n�^>��HFWp�!A�?��\��!K-҆��@�'@�񲧉S�z��b?��G%56����\�u���`�K)��N�w+�VLu�W6�_~��G;iٛ�F�/�o<�k��HS��Aq��r������:_5��C�1�C��u���I�I��Y��S�Au�q$�G��|�\I�Z��%X�"7*4jƟ�ƏM��<�H��u#wt�Q�~R��$̑`����%�k�+>1�b��(�H^���M�8���JZ��O����[�$܉�f���:�L�������}�g�8faa;�Q�Z���rb%�j8�D�(u��B.�HHp5Ӎg�Y���T6��H�0�%#��?R`E�KY��ML���țm�1[�.�9A�5_4�6�{u:p;E���%@�Fk�S0�@Qe0�8c\I�]�9��������4��5���%z*T`�3�����P�K�PNETI�Ǝ~o��d��D�b�g���$�L�Iĸ�!Qj�'E/�m�n��2Ĵ�_������.�(��*�����!�䗹{,�B"m�ݟ��+�:���o�suwk&�1BB�[b�M���&��'���b�%���rR&�����j��:�`�U�}'Y����κ�[qz��F.L �<��ag�������H���f�΋:��1}�60�$�j�=��ܺ���:[��E�3�"B�>Kt���+�^t9�'�72?���(��GQ�FTf�b�0�g�F=5����I�>up�r�}�{s�l3fP�@�&�� �s23kĴ��n4)H�T�G7py"�;Ygq���OZn��W"��A&���1��|`��H��W��0�D1	+�s�d'�Ao��ԝ<�'�F\stE��Y�}�����0�ݳ��b�'�ƌ��d�U�fB�ݞ|͡ZK{�}��!.!b3G�F cK�mtP��x����_3��0b���ˣ�?:�I�f�5�)Xݲ��mȭ�[ƚ���	�6�������o޿��}ô.�%��[Tl3�	��s�b�j�J��o�k�+J�~�FMq"�<�I� ��d�8n�x�'����x�OsM�
�9�.��j|��[�_� �sJ��b�Ң`�`��?����1ͽq��g��':i���Y����u�w�mq*[��X6��;}E�nϘ�}�n��₵售�4\�6G���A�9�2�����]x�=BI�����u����l�]yk��d�U��@�ѩ��#zYґc����z\	{�?�� QHDCA�!�w�ЅI��}���	 ���g+�Y�3��M�t���&�[_P��/�p��W��,�9Hj����C�x���7�3<�e���|pq�����4��`M!�=Xnf�����hqh�"c��E-��v���LL�T��3p:�f�g����7�L�~~
ʕR5m!��7�v��J��O�5��>�}��%����h~�t��]�3DG�ٴ�)��2 z��b`ύ�.�1�����.!z��@�.� Х@i6������T���\��utV6�>�\&Q���2x+xm�dw��e�{�Sl;��3�3�X�6-��s�f���}����ׯf1���-� ��{�*���t�RM��}�k�/��>UͅQS	k��浢Şm�T��ꔓMl�v��KEJ�1�q���I䷃p���ԚZ'���b��1�r�L"��W}L���x�"���E!<kms��T�G�lkSݣ�Nt��_(;Ъhqr�tFz����0��3��6J<.M����<�lQ
�(��rY�zhw�гU�W#�U���A2���}Ӄӵ2J}k��]GM]+I���zڃ�6��֘�3��V#����� Q�."Ui:�.���髿ߪ`<'s���Ld@���Mb�k�C�Wzf���;���.���+ �X��	�vG��}��K~����]�}�����RP��2�?ː�W�]����X��JK�#�2g�E�;������}[1Ru���r"W~}�U��h�CG����������|��]3 h}�Y��_�����6L�+k�1]~t0��X?Q���fC-���ݺ!�W�1t�K�@�=*��[�����6y�_}���!C�����c6ןxB�.ҵ��c�QGu0�bsnx@����M�.@yJ��7���"��-��[i<&�a�R��Y�����_����ϕ���[�=Cv�s��m���kL�p>��Q����to�E+���Ws/Ϟa�`E��nW.7UAfgϰx��˵2�6��G��<;���u�����ƃ��]EoL�>�c�ϥ��^t(���x�1xKi&r��� ��m^2�]er��O�D
+/���n���-{��R@$&?�׍ڛ��Ѭ�VRl���_��좯�+�T�Z:�k�Ϋly6�Ԟ�}n�L�c�����_����]k�#έ{��±!:��n1'��xye�e�59��խ�Z������g}�
�<�����C����Jǵ�/�7-����P����(vh�r���/j���i���S�Ф>�����{�^F�Qv���<ze�����0�v�gi:gH������g�$E�7?m��$Npzi*Ce7�/2i�(֏�w�Ӏ�lJ�5ҽ�s�('��v��1�$r�&������S��tBtR�� S] �h�:���N5��j�$��R֛�j6av]F�(��IY?��^���++Ż7(({��H�B�+���ﴦ�|��p�>�����M��FMi�R�¹������Z{�������"gJДzn9� 䳖��E0� �?~�5$��b�	1��UQ������y�H�ƿ�/�-�"�'q���'G!�މN���M�H(�)�k�3Wuyrw(
����τ��cʢ�rI�M��ak,��V��R�	�s[�Laֹ�EOi�H��jn�
�R�Q��T�l�\|A�����/�aX� �G(\
��E)}�g1�u�/�	�~g���H�Ȁ��[���J+c�"D:
��(q��T:=�p�]���,n�Te{�F:��E�Lf �J�L�Zܹ�1�6�i~2��}�4��F#S�G�'<' o@V/uEX�-qz�T1ek�Uk6	[�|8Q@�U&��~pM��n\�t�����[b�?�ѫ��O:�;M����Z_\B_q�-7�E�W�o"�����=x��J�y��*�9�Q����^�(w������T��b�Ce;���ZB�E�u�}�җ��w�QKE�KI/o�%"ӳ �Ik"���SU>	m�hL��o�-�#���q��[��rFfʺ%t��,a����"Lqߗ�Ow	N��t3�+��Jd��NKi�T@'W���yk8���wZ!�G�ˆ5\|W���͈!�f�����zԭ08�u��d��rPD���X�3�c�a�YHĆjt
3��٩O �>\� h�WXC>�-q=�$!�0C�|Lr3��� ֋�eH�?���8�:>	��,ߞE]�K=�t�ɼ�ڸɺ���������Hf�h�Vs�\���J8�8�ǐ��'�;C+e�oU�yz\�|���,��(\����g���$l.b�xZ7��wG��KB�f�a��)}l� ��=�SZ�f�DJ��靊��X<G�F �������*�rn?��&���Q�&ōuT�Gh{����P�ca��X$��+g�`v���#�%�-w����.]PM�LY�C�k��S×;�,�� $��44���q���r3��\ �v(J̵�oaj���f�:�r[����6���{�\�0Cj	���0��rj��[>�ߥuU�'�w'4p��C9��r���g�KtfA���	�i
�#��o���>klV5F�;�S$��,	�9�@QH�Ťy꾑��VǦ9�� �;q�t��Bg��zasƼ�Of���R>�k@+����iDihFCo6��)'OzaOh��D!�z�Ε6t�lR�
ϯ�8�;�E� 4X{�1U�g��QF(�\1�G�#�Uu�5�m��dS���q�Eut#��8rh��q�81��y�#{u��uS���PN~js��"{C��b��	*�alM?Q��ў�TT�����ѥ����K/e����+�������m���0iz�}�Ƶ����q[iD�C�㻻+'�]f�Tn�9��'ep+m�^�����l��|�,EfR��ԣ�l}iԏV�\:����Ώ[��EbK�ێ�g�5�ʅ���q�f%U���x��kc�A�{ʳ�LL��ϯP���j-TƎ�5A��S����Z�A���M��{���;�Ry
8/��VI�O?u:Ѵ��:s����=)T�d���� ���7.�x y� R��Z^hFat�d��9�@lk�y���G�1�4���ϑm�3�(Wz�����l������Q��i.�[��ݑ��p?�#��f8�����ָ� �A����<��m*5�>�ѷc��v����*�&<�$'u$�����K����#��2�v{zE��L�#Ѭh�9�P_Ez�J�=-Q���wh��g6��2[�4��U�fO��&�5��Ziv�lk��x����;�N��L R���
�����)���Jz����i=RAD����/����g�4R�%b�K����F2ojE?ȟ��|W�񠾨���6�I��*�*%F�8�8�F��Cl�̆�+����n�(��v?�����ۤ`�oک;��j��n��a�ܙzj���j�g��G�B�1lҙ�eڽ*I���(����)E�}������N�ѵ�^�iY�������:Ov�w�ُ:���j�M��}X>uS�b,VSQʔDo4��Gl��s�*�l�"m�C=��o������?l��������Y�uo*p������+�f����3dߖ#y�A�kǶ��L�����93[qs�Oo	�hG�3J�0�_���`؇��S��P�HӨ
�^1}'d:���9Ҋ �®!������$"����R�D���èS�K��Ͻj���C��家�
r�������+V[�7b@Q�8���1�Z�R e뫬{�����(�[�+~�f�t�{�������d	���N��">J���1�
���]�7w/B��g�zX#����~WH�2�z�V`6�mk!Zʋ�>p��7⶟���`���P�m��2{�{�j�
�(��Zw!	�	�)�H>=
=��S.o`����gH]HU$r:&1Z ��l�2�U�xg=j!B|f��铤q�x��N�LJA<g]s"Aٿ��W�sh"?�&c�-��,�rDL<A��c���^��$Ļ�W9�i7H��ߒ���|��Y�vm^�|� �0��%�Ӫ�1�l �"��R+n1�&�A�p���Ia�T�1/\x��Q(��63�F�9�,K�$�J�5a:��b��}���0>������+0�G��Z������nw�K�f�W:�c�F1��W�
�ϧ����m8i;Й�c�r��r��nw��P��-�?=��E'�<��Am�h/ď���0�p������x�[Q}���)�#�L�oh��R���)��N���b��gˊ�L:7�؜����_n�<xM��>~S�_��gb��l��c*,�y"��Ieއ&|IOB��Cs'�W9��	m(k�V�\Q]�4�d'E����.�s��2I���%dSu%���VEl��qm^�*@���X�	W}ͨ�K�[O��y��ϊ��ڏŚ�!���+K�2������մ�>"���,&[hjg��Q�$������<>�MqUX���0��$>�O��nPy��Փ#MCf?Gxg며�d�A��Q��~$�d;��V�� .�Jdʑֈ�����֨O�aĔmv�$��)!���W�4�@���ו�iE�L�6��a�-��|�\�W�.��Fs��ֻ��U鍿&\�D#�g���p��Q�CD�aKC��� �q֥|��7��`!@�S��O�Q���l�c��:��<AQO��m�HX��8�7w2E���Z,vK.vd3'�Ht2 C*�Ah���i
�����bB��Y�4������Lj��lou�����Xu�%/��j��&�U/Z@�r�NQ�Y-��Fz��NK�R1G��z�㧈U:��4=���&��%��pM�Ba8����E����m⩓��@��@掣�e��5*����b����
y1ee�E�D�JgH�vj�N�i~��<�T��@�	����nk�^��ڗ��M����y)cO6ǋR��/.s��(wJ��}�^�6~'#��`a0��:�Id�X�ǰ9�{+zG�x@E�#?�E�=-2�j�7Y����^�����]9�_�|Q�q�@��,u���kC\�k��6�K�v1'K��^� ;��]�;}�Is��g�xv�/�I�;���\���׼�\�����&�j���j�*cX�^D��(��;�c�d�h�E���W=��8�M��>y����_NS(r�J̀�],?�Ց����u�ln%·'�6�Obt0�Xhᚥ?y�`N`��j%ͫ3��Ӻ��P�1��Y�I�Y�*�����+
���szc���%�y���x�U��.(kοG�6(W�?U>��e���(�tu2s��冩i��M�m]�d��K�_kȬ�:,g��X9������T{�¶�nr�3#������A�չe����H���e��EE�\[pce�:��I��͆<��;����/��.�<gطת���ed�_x}f4������{��ESaI�lg�0�\y\��w���a���(ɔ�;�}51��/�������*.��q�Vv×z�#����+���|�^�	p��)��P�WT�XO��?3��{����$,e$���[}��D;^1�C-mp�����vF�V��5��	��|��[�D�Ǳ��u-7&!��)�v��C� {���2ׄIt녻'���~��-�����2��Å�ch�6O�{�:d���='&o�.��ۯ��y��h��A���9�~E�;��~���7���L���f�	�U=5�m�E�4�r�km���R���v� ��r�)4{궝�oƀ�f�{������Q�[�a�q���E��j��!eREj�b�y\�奞,��9�������\ ���o����kCċ�QE	{���kC���ߝ�ՠ�����~D�.j�K�u����%�Ɛ1�_���.��d�-�>΁�����{�)<0q�r4y�5"y�<Q��[���+�&؞;��t��P�ӈ�Ź�&s]O�	cx��4u�ȭZ2����'�ܞ0A/G9|�S��Oi}����"p~�d��gZ+��"�y
)��/#.J{�J��Ճ4�~̞4_������w�i���%lzD����b���r8��:�뾶`nB�L �`p�#�1`�#����M(�!��m�����m���F��`V#S�������,0��P"���s�en��f�P!���PP?cd,�}�������{��1/>��L��N(ņ��K����Qcژx�n۬,*�،��V�ߝg�]WZ?nT��;����À#�,o��˘�������#�ٻbȍ$�̗<�8՝�A���V�|g����z?k��g(C�������kN�x�#cD���X�M�v�5�3)�Fu��;]�<��k
����C���I>��U�6G�9����ІǊ��|E�\�Uy�XO�{7g�S`�*q��L����c�c��������<�P{��<��-52SN�Uaq����upW#ڊVYhS��\Wzu�#����Y�d��.aW��h�N41�"����U(�=Ӣ�i+���.���֏ ���@-�M���#`�� w,Uyc�J4�F  ٖZ��>�K��^�{"tV���@���V F�Bgf�b�˒��s�f�H��Kߠ^|^̕b��Ј���09�Lf��2�a����'���i(�C�2e=A�g�����Rg�v��lH�g�w	M�I�M�;�ۓ���A
���<���'���{�
�g�s�&��Qs�1�X���`4 (z�C��,cCu�(������-�桖[���$��'yLiּ��q�mM���U�;Ԥ�g�t�f�c��+�{g��l�9n����:'�)���E�S��G�����H�蚫}Lh(	\�w��:6"�����K|	�������]��t��1z�������s*���>Jj�fV��&:���<�F���oz舉��v-`f[�(8����ү�ʠ�#�Qi� BLu�kۇ��e��W�l����{Y*V�o��4{���ޑ+�Ne<z-���j�H ���1��[��.�wIw�X��-�<�d�y����y{4��|�I�._��S݇@�w_�\4�@�8�C#�c����d�:�d�b��Ep�%����hƄno�I{�:pm0:�0
VG
`D�J͍Jc:�f��rP�p�p�CQN��n1������i�:�	����X,�J�#$�����XR^g#a���<�hz�+Yvly���� b�oo^�vHn�hpn��Hxv�\e����N����'�M���
� �=�p���τ �n��u�5�V�&h�׈>K�V�H6K�5YRRҌ��U�Jy ån��$n6TD3$�D9���$�J�-�p��H�Ȃ�W����UC�������=_je�^��>19��C���uV�V+�^���E���ӛ��Z��l#"$_� U���C���0���#��Ǵ3(�Z���R|�PÊcٓ�;n2�N����k��f@����$6�9��'I�+(��>Η.��K=�#5I�e�yu���t@Y��w.'H,BIl\���-�֪I��^8��
���M�=��r���v�19��wly��C������A�M�f5�m���?�)�#T�0B��qm'[����娝0q�m���I�O	f--�!���	���Ѫ�j�x�t�q~kr*�~��|�!�6j|	�CQG�7eC�5� '"����L��}�����o����S��G��c�n�v��jϮM8M7�rV��bI�qZBgt���(�QQC�OP��<D_���|JY��4�L9JMc��:��;���q���¶�XM���\�x��pF�i���-'�	��Fou+g ���<��u#+Ae��,��i��Q	S�z��ܳD�������BW�N>¬f��9���^�H���_wþ�0�����kz�]�� ����{�y�z��(HZ��dY]VHau�{��Q���QL\�M�8 �j�aٱ:�K�������	�'57��=᥃PV��T�����w�Q���3�����D�=���2=��_�HKގp�D�!x�t}\0B��&�gǮ��7�g�lQ��-m�f�A6ҏ\��dgQw��qyku�7�泖 �/V 6�۝~������@=Erk�Pʮ�"�G]�)"`��C�ϐ*��IJd����%��ּ�>����6LB(7<$>A�z�s��v�K���3��1�erV���%N���y6AY�hm��NT2O.���:��2D�{�i��&�������S�m�L콛'����d�dk�w�L�K���ը��dBY��L���da��e�U�NWK[��ޅ�f�w���+k`���W��	vf�腸��CK
6'8*�&a�L �3ȩ Ѵʪ�N�S+i1�u�*���n���o�80�� ��ͻg�C��s�d��
lL��fp;V��#�IX ����j�^�(2Lh��4�$g%�MND�'i�rVl�?4@fޕFp ��[c�̺�[�q�q11-��~�8�k2l���#{-F��ºF ��M�
ɚ�#ӯ��ŞG�db����u��
����l�����mV=�Q���|K�d"ӁBꏁ��w�Y�+ik�4��8h�%V@5���g�����"P;�c\�D��t�:��jcu�ݬ�<U��:ީ݀�R&�wvbv�i5:�'@S;����j2cp{m��X���zM!x�6�����-x���2�v{��@����E���@�"a�!�����!� NJ"P�e0~���3{���ݤd�t����n��򰙏�z��&�e�Ɣ��|�'y*18���5<p]˂llԤ�}"�ўR����\���A���Lx.GnKB-R2��jȉ\��`Q�zX�F*�Gd*.
N�XB9�Vō^.W�/7S�Ho��aL� $��)�lw��~�-s���> n��w�⿫��Mq-��5�R�=�Bi��w`�ޔ!tG����7�4 M`���bu�J`l�;m�ŖvJ�3[)��|�м���=X�n��@�\8)7P��;�QҪV��зHn�I���.�y	q](@o�.Σ:�Z���^[t�2��EF����<j�Q4,�y��'d#�B���ۙ�$�������z8ף�,� 1Օ ������]�Ń�^��p�'ܑ3K��I���$�7.)�e�:��Y��8��s��7�ڈmj5���a���r8A�2mۨ���ľݻ�.�9i�r� ���]��]m������k�҄����k@w���(ro�xw�&�B��S�������@ �湱	V 2��mK����>�o�5W$���6M��60���hh%�*�s�_��b�-*_�T領��X����3���ۄ�Y����h[q��dviJ��p=%Ĕ��&0q{��3�~�(�����ov�4�Qнk�V�/���Ӑ���x�oGji��x]�Hտ1��xN�q�x�a�\U��Z�H63j�|��~��f�v�
ڈ��&�bf�ȟ#t]��i~��IEG#lUA�޳Y�����R-&�r����=ӗ,��Z�Wp�4sKU�ܸ ��R�b^��^'�T��@��`�������j��BLuP��|��GgTI�����x��@7%�h��窑���������m��w�P4�Ԟ��O���G��J��2��i�[?��8_�h�H�kc���ԫ
LE�ռ��R.M�V#@
�������P�I�=M�l�D��[�*1�(���Abgǘr���=�+˗@Z���e�͢��"E3�×�����?��F�̙AYU ��`l	V(�3N��1Y#�8[�vs�#f��쿸c��Auكi9$�j4;���u��	���}���Zh�o1�&+�9����#����t��@�E�xK�8뛅�h��z�jU�l����X�0�ע`��r�|k��E(}����#Җb��r�C������� L0�$j��_�%a�j�A�Ix���� �t��~�;��X{qCF;���Y.zt��OĤbw�h��z�,� �l���=�d���8�3D�����|=k��Dl�b���,c�<�?���\=armn-�;'�7@�*�M��s�v�r��4DR��$���`q�K��� ���D؀�]��ͻP���2&�R_U̙�$W�0��A!��cF��)�ނ�(-Y�N�Z/��wru���~����yJB�������Θp�Lh=9�ʺa(����`�F;�qPqY��n�j}�0��WGk�����A�)E-�Ri�B�W��A�cF'�"�Tm�t���{[e*�Yu[p
?%�(1q^&����-x��+�}Ze��CVj���^���mG����n9��ټO 	&n�P%[�G���w�Ծޑ�.i@qo�˻O�&��z�#oaKc*M���DO�K`�/��Y��5F�Ԥ��=~�~�R�Ɍ��C�����3p�Ì/��r��Y�*̲:�b܂�H>XiK{��4.��P�Wd�*�j ��]���$8}(�q�a�{9����M�+���
VN>�u@:/BR)i�<��Ȩ�e�gdC�4($��[�	�l0��/���Qw�������9��@�[<̻{3��Bm���������r��O?����Y� m�t�["Rs��-�-%c�Uz!�=3�@�'�~_n�|p0AG6F������z@%"�C��MrRK�ף�"�E�m���o/�[�肗,}���؈w���"὚�6�$����.�$B�p�5�z�Y�������QQO;!�)��/�ǖ������N�Fk,�O�|��%U�c+>llh��׮�$�y��lZ�e����U��?�:��������-��7PW�%䵴9�U,ݭDn��o{��tN���MV�wk����k�����?�>'���)���Z<��r�?]G)�@A�%q!P��?�u
��f
s�u�����;{a}�W� ����P��M�q'��.P�Υ����Lwkyg�OL�>>��� M�p#�����*��7�(��bZ�e���Z Ք�5��*�i�MJkq	^��4
�b��Γ��3̐���zķXO����"�;(ʢB����h����:�������(���T')ё+N2��q�Ԛ�ݔ~���^\�����t>Y	����gr�S���V���S��p^�!Ț7�Mw}l>~���N��L�p��P)����V�j@"�ΘE B����μ-���f����.�B3��],�gA��T珸�������f�
�������u�tT0M ��yi�����_����z�Tso%����E�rl�3�2��G�Ӫ^ݹ�>W�E)]C�E�3�t�++�	��菉�!��{�)���r�gD�ZxPc�����o��L�jc�wX��Km��ǯ�y�͐#ooX�������[C �`h/�R&ej`�$J�KR����1��3�{�v]�FS($Np^$l����сnB.��m-4Һ���c�m�Q�Y�ʊ�D���v+�u���m�4ˌcŅ��S��UQ��l#�/��.��X\� <@';�4D�,���O�9��Y�Ze�C�y�����X�qޞ0tL2��q�EB�z���u�,aO"���-��I� �Ae��B�C����� bw�i�@T&c���^��>�rggW7or4�!���h�M+����d8Э�S�D��T��GEF<}f�%�7Q��ٻ�H�vX��Ŧ^:��g��#�J�c������e��ꊚ���6���S�b��sm_?�8U"ٜzPB_c�&�]�P�>�����C[#�yP�W��M`t�H��|�H�}ىz�BR|im<klO�klÛB�pΑ���R6������N��B�t	3AT�^��@V[�3�8&_��Ť��#oZ���hN�X�l����|T�~ąnzm����h7��pg��B�/���: u�+�kGh�%��+E�[�Y��͛�v���w54���>�}���o�������jG����°S�M؎�՞�|<���vl'�<�g�P,2CsG�O��؝�"��G��4 v�e�� c��	�\蚌���:1�ö����Z��wt�f���rŎ.�.�=��o���'�\pE��_H\E�f4�#��I2�yU�6e �|lb";�`]�u��� |E�h����{�RT�y>G�:�7��54�-���j�M^�)���
����Q~:���'��ۦq��9�䑧?v��؁S�tt]p̍�më	��uwE�^�[���R��X�b����P���TY_X����oж��p�M%���h9��'(o�#[���e��~�;6�������U��6�=��G��P�t
Ҋ	s�5@)�j9�W���!�ʟ�X���^�V�Vɭx#�<�����?h!��T�����K5ue��zJH����F�aΓ�����BZ����<�&����Ŵ�c[�_�.=<?�r��u�#}웱X�E����K�'[ӕh��b 5�kY�s�f��cY-Byh���A�ny-MƮ�p裧Λ��u���G|}Y\�׬���Q?�l�jr�S!Z8��ODZ�ө�Q��%9����:�V�����aq�?&s:΄W��G�~ScB$���E�)le+���@�9�S??�M����Eբ��X7�@�I݃.uz0!)jpҚ�,�jq�0��e��@�M:�>	e?x"'o�d�H䢕%��`���ǲ�n�����"�Tz�rj�f�1��-0��qe�ܡ����A�N|cѳ"����#��E:�TP����e�;���E��E�sӃ4	:��@)-l�(��,�qN�9�!��D��1Wllw�M�!PJ�^JpY�e���e��>W�I|��z�!?0 *\/�8�(�%���,��v2q��������>�@,jwb���ܮ �9���n��c��Y�h��4������~@I�nzŸ���\��N���dɛ��E޵�&�l.�M�x@<+!|p�S��}� i��������瘈��0���w�����o�^�A���!9��i|未~��)�~�NA-��+���IR�z���I��=�U)W�ǻi�!��	]�����,W�hn�[�bz+�M�����!���������Y���r,U����� [�����r�}1B��޺�$Ibx`�<w䂪���R2�?^�O��m�u^�.�zP��`��ѝ��#W���ܮ|Ty[�n0Ydm�LZc(��5'�>H��7rDQ̀rf���a/��b����R��ø
�%4^��l�p��K����s�Ŗ�7q;�F �3���B-f���x	���|��K[~��"I`*D�&�P40MO���LU�9������2 �
�!z�v��PG-��{r�P6��=W#K���X���R�b�3��C'x�r3Oq'�b��o�y�5~,��=��5�]}�ߌ�oG�C���PP�ll����A�� `�BL)TT���5��P�ˣ2kY��������C[	WS���koT�~����d�7�l�:Y $�A8n�7_6Ώ_�8Gi�ݗ�0���������Q�<�raе)���jK�_/iy�,�m$���s���Fyd����zǘ@QE�U+�B��Qu|�d�fZ���X�'� 5$쵾�Ƞ��>��;Z~��8;�/����0�:�~�,�9ۑ�U����������_#�:CaN��}�lL���$u:��Tx Ȼ����n+悷�5#m��[�U�������(�Z��m'���ܶь���i/���qv��S�[�V�&����u�C��K,IA�R���/�3p4GdQj��+�1J�e��gn��ׇ��ĺǴ���Āh���UD�q2\}�nq�ˀiUʿDE��q�ZcH<v�wM����C$��}`O�B�1�ԶCt�[c5:���_Ix�m�S���jU��˜[>>�y���,qc�FH�9[�o�>�"N�6�c7ř0��v��֤^b��)�P1����-�H��[[Cc3�Qn���ל��m��Ѧes����q���n���"'��_E"-Z��q��S]��\��l�.-F��1A5���I�Ѩ�@lqp�r��/8���W��dW��"�RO��_�J�A�c��B�G[R��K�M��2R�0���A�Ű����`��(���'o�#:���ݡ���t���A*�5��I,!�ܴ�[	������#z%�0o`9#�=0��q���mn�6 G��f�ҩ;.��?=Y���#�M��=���Z�/�ȸI�T2��:J���}��m���K�P��%��V��}���M�QwC�B��B��k'N� �����R����1���O�0i�J��t廿��Ij�-"3���J�vN
��^u�,Gr�s�`�����O����u⾋�W��#B��وq���#o��v�R��ʉČ�W��ʴHE�1��S������Έ�XH�-���!�6�'���R()�âbޖ��fx}�M;��@��5[O�&�іЈan��z�U�G�ڄ��۸Rz震ȱ���f���wkv̈����+m���Qlu`VFvB(�@�S�ҁiG�M	PPrD�]��{X�V�z>}*��t�!;�������R�����N�*Q7������Eµ;po`�nr��Q��%������e��\/"�f�����F��/WtycR��Y�O�u3�dO�+P/{��&�SW��أ��؊�N��а�>��$��b�zK����!�w�DL��.8�=����3FK
�e�Q��I(!Ѻ0��$�wA"��b��v��;Q��zAl5�ݚcȇ�j-����l�� �	���$��I#��e���D��p����i�YQ'�nD6FQ�Ǳ%*	6Է9�Vz�VB���(d��5�-�q��(W�3�u��&ߥ��&9�Mh+Rd�*��6w�#�i�R�FF���3�ht�0��R���d���t,�`��I+�4�ƶtB�'��M5����ր��:[�yMX&ʯ$�x�p2�wRw�UM�&�Ӷ�O�W��e/'-]�D��%�A׼�G�4����m@�0�-1xD�#G/�2���Z�ޭN��O
�Dhr��쾩<q��q�O�D�N\���N��h�kƒ��4�@��E?��
��w���,J��p ki��\A��``�:�7��a%A4O%I #󽯶ľ�ꎚː3*������NY����=�'�2L���4��q�[��r��ؤxAAV�_L�m�؃W:Y���N�:�T1M�t��5
~�W�*ZLk���N�U�PQ��G�����f���)z��I��,�$�z��k��~�d�����2/8��I)P��ܹ5!"-�up>Y�?�M���wr�#B�i9��m�۰:�81n��n���}#��h2{���޽����4<r3ҧ��,��<vk?���>k�@3+�qg��Pg�,�Ĳv�O��g*/�	ni|��pki"�'JG��
3z��+��"su�P%O� ! �,g�����Ӎv�mv��ú|뎧�5|`sG̾�0�q����+��� '��ߏ�-7[l6�@��_p��bgdf�����)�o.<(�(��es;��\5�ࣧC�lM��;2x4-6�v���s6�����?Y�'�n���֣{����O���w���2w*���H��>��SSKt|-��m8hi+3�w����n$i�a�}IÉ�]�j�r� ����v~�ٳA��q��'K��/i)�.�S�ˬf_�
�E*Á��ǮUKk��s�#����A�֕&p�MO>��!*y/a]�W�j�<Χ,P`,�{j�^}��:KK+;ʘo�1���X�Cd�^�Q�1�o�w�r�S;�',���p�,M�ze��'���" ��Y���%([��<j4_%�~K%���찹*�<&sG���.������B��j��ⴕ! h���C����S ��� ���~��c�d�L��/+l
j��A2GU\L��󒉚x�4)>-���H�o�7:�N%(F�����hA__��ʥ(�r�C'�Z4q��\��?�&��s��_ ���̇^�)����MvQ��u���c E3�$Po��.�p� �hJ��I.i�?�u�٠$�`@����Q�^�Z>s�)��;��b�Bø]e�VS������6a��lw�Bs{̹4���U��4�p�0XdcikN>C[��WZ9�I �<��+�=��B�' 7��<�zL5�Py(t�������9�J0�����4Ii�X�s�Œ�T������&=����f�AD��4}AGb�L�LT<�~��{�*�����#�_����5Z���cc�� =g��(o�m|��-�χ��A�/���g�w���ze��BjkA�dV/W��g�V�0��IR$+�B]qj�W�`�QnA]�;�+� 7V��F��mg�j{��7����](��aO��rƲ����}�c�n����RӔ��Ю���WG���W�~�����M��I�U��f���_�X�_���-�>p���LX��Z'M�Z�xW���"E��d�G��O<���D�;�����
�m7m#p�cKt E-�G�_�Е��Ofg�&oT��ㆫE��mwo:l�
�B'�����w{�����_���Y?
C��[g��9�y^�1@�BO�ר�;���դ?���OI���1jbث�����H�m��''!Jh�~Ptڏ��nx��m�����"3�z&v�UWnL���>^G^E��>.0�*��"��ј惕䈫_6S-�u�M��������A]���]��n����	��F���s��,vI�N��Ͽ�D�q����i� dw:Q�	�y�h��3��	��+$�#�ɘCF�H�FQ��Ms�a��Y��c�B�HV���qj(�#{�S�U]���_\F�5��z]�U��3�JK���jo�W?~Vy��~%S�da�3��~j�%)��,�g��~�V7�W��(��fm��:Γ.�BC�n�͕��{1�h�2�[Z���l������' ����u��7�O�����R!�?n��PX�\�E��hQ@���`m���Y�?��ġ�EPq$E������ŬD�lL��i��W�u	A�|����hm���z�A��}��'b�E����b)�-�^4��B�ebK�z[R�'ES�0���������h�����;æ?�b=r����m��J鄃��ݝ� ����5��ݽ�k$	���/�L�v�J:��n� ӫ6��푸����8�����^��+|����]\80�;�=n �;�s��hv2�nvZS�}�>[��4w���x'°�/�����Uw�=
�\4��ޣ���Xw0��V���F(��[2%����6~O�0N�	�G�������<�gq	ѷ9E)-�\�3��d�쪥0�Z�W�w�j���$�r]�i��E�R�H����]7�|!׺`�$��s3)d+�/̾w����u+L[� qۡ�_�����m��7@y�[R(��橶���s���p��5Φ����߆*ߢ�_���]n��m'��ng/��!��XOg���kY�a���px�}���X�g�����,U}��IҚ2���H��T��������8ꖺ]#��ޝC!�	��o�N!�w��7�Z�7S��f8����E�=��ۤr2tG����IXqd���� 5� ��hI0�����o*D"r�ţ��9Hy�qrX*9�H$w�Y�aKy܉Ё�����w|G�m6���Qx�X���^SiH�mP�(UI�Ws3��J>�_�0�;�P��H�0�S����a^I;4�.��ӃB��\[jv�:vQ��`J����]�ه�L �u?��������GH�~�myo$�Xh���l�<��i:���H��m�%��ڝ&����}ʵH߾��v#V��="}��;#g����b�z�����[�ڃA��b����W���3p�H13e!�����.AVw�7A�_��%t��w��Պ� w��xf�K��k�:��i�dg�)�V*�뛠���	EA-F��v9P���I��C��F�_	{��K�eB��o��QV�P����}~��nzݙ��Z�1�,���3���m�`�3v�*�/�(W(8�y`��I^z4����v�piOE�����#+>��(Ĥ��i'AH��n	�/#�j-J��+��j�)�"�݂j��c~?5�"!�o-�=��q�uǆ�;QB�� ��B��M��u���S��$����v���)15��e�B^��yA,M �|,�ٽV��_�O&�G�Qxj	�1�r2!����쑦��n��ia�zx 1��|=��>����K��*mi�i�K�RSNc��;+˾�S$�1��K	%�=�?a_A�B��wj3�X?��d�l(�?�K6��iCKR��$�ޟm�.�W��$���GCBU������ƶp��^ML#�'6�б���&҃)S�Az��oc�n��k_瑐�#������K�Rx$��<^�+fM�2��T���=��� }u9�	$1B���X�;Q���gQ��-��%"-��m7�$DX��yʑ�p��^-�u���W���ʫ��_����;����E�9Q���ԅ*Z�W-}:˾�sal��c9����dtM��C��Z��IF�7j���=�5L�E��"{\Ω�:a_Lެ��\�[(G�o�n��ߥ��.1E�x	 a���5ŚzN��1������"a������a�e:z�Px@.��(��n]��e_Q�񷫌��2�h�����B�`ꑅ OK*e�m������ԋ��1�s,cp'�W،��`l�T`�/O2{*�o`ѹn���s��\�&�<cnز&P̀��Y��w����'�(S�r�D�R[��$X��/Ope�To�|�E]�К�����f�*�d���7�R���"u}��S�C�vk�ք����Jjh��4D��W5�8�,���� ����b�-�-7����,س�i7^�8�</
�}�i�S�BM2�_�,KfҪ(�m��k���_���n����~�ۛ*����6k�1��̰c�8kV*��:s:��.[pkT�₷��Ǌ��$'�m��iz�a�I�8�xw�s������g�n��kYD�>��{�8�!S�P�����o��!�/�V��AC�ֵ�+��Ǧc]�hҦ��r�[�zz��ؽ��M��J�WW���^�e��!Qn�v�p�O�����r�E��L;+��\e
��b��_�jj�$�}��G!�����F��m�M�q�M'o���S����"�O��K`��p\���u�H��Zo�̳�$I��+Kcˠ�O�k�K���U�7!�?���{��[]���h! ��&�Q�q��-��%���RB~�� ��I�d�s׵�w���JՓ*Vl_=���j/~����E`e���x��˶iI3����.��L�y�N$ �1�����+R�s�t\����v�
JV_l�����{�F%�����Sq����0r\p��O�b���uh0��7����͠x=n��ͩ�[�����R��l�\X��	m�O:0�QM:���GŦ���e�'���=ĭ��1Y->�פ��T(�����<��rA����Raŵ�bP.͈�6�WH$U�̣Hz���7ˢ3#nޯq~B>mZ�2��Ψ�����8H<e��]���O�:`S����5KC�U���e֓��PҌ�2���SLl0��].�x"�n�/<|��?�j�zcU��D�P���hD��Κ�;M;0�?�l(lux�r�tn�&�8����w$!�^Y��{���u2�E�+���t�'�__N�3�����spk�����y%��|�H��[��{i� YuOĖ���T���տl��f�c���ڌ&��Еm���?���%�ġ騔E��I�ϻR~��#�|d/�sȺe4�� ������+R���������Q
�q[�z�i�x9������v]�Dn(p�X�a-HK&��)N������y��j_]���k}�dN|��T	�_����ظ�
�lW_�$IA�Bp��������i��r:4�i�����B�2_�VU
_5ѹ�!�����Y��������T�Eʵ����՚��:��������̵�Ss�U��*s��@3��=s!c�@<v�"�`�,5����HB�!(�>`�0�I(�%}����F�0W�T���\�NFN���A�o1�[4�3��Q'�%q���]�V�5�h�H�G�+��C^\�W1�C��f����`聰�{A�$<�c>|��M6��d�����T>��t�U��=* �������*��kcrj��`�[~��.̆����pC�<�9�{8!Ei(���Ld��Q[�N  j�w�AM�?հ?���ŭm�)�R�R�)e�s�>���:��nh���s��8�F���N����Y�)�©k`��g|-p�,W9�Sb�%�{`=#�։L����<�����o+�$%vU��j>)~C �Y�bJ��=�4����ǜG&���7dA�+��v��-5 fx��Vq/�2��e�}�~���M7�m��9R�7���t%��\vh{���c���gpe��z*�L|�*n�V�v�e�):�l�����������J_��>�ku���Q�M�@����Ās5�C���Q�3�OmZ��rZ��% g",�(5m:����&zDH��i�T��E���	�,L))v�T�3u�b�f�n��R�Աs5��5��\̺@5x�
ǡ���#�Yc���!*c���@T^v�H zWkTY��k�#9��J��ۤAW��5�U92j��X؞HL�pޜ�6��|Q�<�&G�7�-|o��j}.6���wDw��*�+c�(�z��ɧ-`��{*��.��B�t�|��THf�~�OG��?!�.�dk���r��$�H������ì��r����0����A�QD�` *8��7�؉�.`�$���@�2|���w��T	2~O�z{�H|	�k����Fqf-��/�w�8$ܗDv���k��~���C	X�;�_�uk���n����F�����l8C�9T��~)|O܍���ٙ�K��%�f�Ԍ�a�ɼ*�\�?�oH��@�E3��N�b\b��<½z�\�P����"�k��Znd [7<�� � 6�a�4͍�#/�w��a�����<���͑!S�{3��g-z�W5��l�6q�d��<3�9G��x~�	[H/Y}k���1A�*	ƃ~������@�*�<��,��1�#X-
�UJʖ&��#���z�B^�,) ��nUn��`c0ꩢ.��IG�O�>V<���M��ˏ7-�C��$�E�3���+�L�N��K��ie��1iT/���:���Y�HO#�ќ����\(�C�1��M|(�����i�K����*e�`��$�7çq�!�Gn3����-�~koa�ڂ��?l��|��Ƹ���h"A��Em�8���2��'�1��ݺ����U�������M��D�sC� o�x.Ӱ��"C([��vTњ;�z����*>���? ^�)]u�e�t�'ҝg{8�O��W5�TL�
�C��
�x:@;�G�i �>{�-W�(F8/0�7iy{1���K���`��8���1�ى8ĉw4 �V�^$��C܈�b�?G]���7cUg�<��Įnao���W�=��O�k����˸ǋw�d=~�`��V�|g>��_�CB������BT���Y��[.��UJ�YC��;@@���-��1�nu-�U�jSZ�ܜ��=�0��O��S}K�aL���n�������0k u������S�Yq����#����ۍ(�<q�>(�!$)]o��s�8&�����s�Ƅ�/�ǱE�,T�WsL�9�ΒV��o��f�L^����"�3n-�"��9b�V����wM��!�Ta- f���J��,L��̚p` �C���M\���U�}��V�����\YL8*�����G����{�Ð�Z:�-����A��9Rn:�@��o�9i�wzLu����G��R?͊���*���:Ov��$)-멜�;� 5�ڹA��S�:21�����Bt�3Q����G���&��A3�ͽX\<�� C"{Z;;�]�>R�-+��$�Ir%� 1�����ϼ7ya����34��w3�5�e����&�ϦdXw�)*~�J-[�A͋��l����];�m�<�{��{#?S�.դ��\6	�%LT���cz7����q�o\��M��Ԫ"ja�c$xN7n�&�q������ۓC�o)=����h �� ~J�ͽ����#�FY��uJ )F��*�P>a��9$\��c�5Qi4���L?A�G{ҥ���Fs�F[�[�n}XCR��~O-߶��~�D&���{u{���d����|?$d��K�{��Q+<SUv�D�0Nx�z�h����P�e�θ�t��=$���GRg�'GAl���}���Zc�,�|s�BuN���Ց�����_=0J����g���_!T�z�<dB��^�r�����#^��o��1)� ��0����s?�+���Pm�|��s?zQo
���9t����^ˮ��p�V���bIE��E3h� ���Zx�@8�#POl����|=�3������z��;:Jx1�/�0�V�(�r.lq.j����n]������g���Ͻ�-s��DN�n�<c��Mص\����<�d� ҕ	,����%��C��E�]@<��T�>�p���ԁ)��d�n�ɈVPڑ��nŷw��/Ci����� =���������i�ÿ���Vj�7w�=�����f	��HU*�sKش�p]C0����n�ڠ�q'p��$�+����L?�����FĖ�bVK�"�>P�W̯��l~���E���fv����6 Jvb󑓃Iۿ=�}��h㥓,�M2�41 �fU-_'�v��h�- �&���� �ޅ���P��N�qb�f[jb�̋�F��'����F�Mh�u��x�ݯho��h�[�St_������)^IUKn��y�m�V��(̔jå�fRg&>A~Zf�׉��"�1��y�5���k�C'=*�v�4i{9��D{$c]1-��"�\��]Lk�}���`9�K��R���8GK�R�:s<�CM�F��4#�~����c&%� �M�:pW.�&}(?�-��m�)�ROoQ���V����h�����>������w-\�E��с>+q6���_��i�vNAu!�\��X��8��P9����9hv`݉�G��)����ș�E(S�����w�e�F:�����K��rW�7ꤙ(7!��q�J���ƶ����v��$�|wAKI~��>|�JCB+�9���+1&�ս��5���̒�ˉ�$L�����α�CD��b8A��"t�?;&M�gt
�Wi�͉U%�l{d���nv�я����t�`��Ú�2��gC��P�!p���&%H��˙�H\�����'�.;2��KQU漆��/����F��ij�T^3�&g:N��RP��d��o����/�k��`x.��'���[�SwJ�	ۏK��2��p��	#V�t��1���5���gfT����
:v%��Cs��2X�2�-k�"s�[aꫝ��'�i���U\-��*Eq-��3��w���h`���Dn��f��'�:�u�;i�R1%Ӆ�AX���`��$	�J]z4z��/�*����+^��M =�ŏ��A�b{�$ԁ2H������_�Z��GK���8��Ю	h�<�J�{ ���`V��j��k�;�t�O��\���C���:���#QW��.��c6��-r����+��ޱ����[����k1"��d삘xa�&��d�����엚��K~n*�%�U�C�n^؇I�_o����F��!���A�Ye�0H�b�ڗ���+97����� %�ۼ�^��߳�F0NC_�+vᷩ�U=��;8���lt �)�}3�t9[�3zpi�=�D2��Wݠ�_9�њ�#H��
�`��+�C�N��Z X1��K� �\�Ұ1sX�?Vm�:*�XrBXc�#���Y�8��`���f�%���Ļ]���5���+��e����i��-"��+ͮ)�����v�%ti���`ZYQ�k�H��e�����lֻ~Y�!rw�@�~t�%�IݰE�ڸ��Q��������n��Mc�K$����0����Po�"��.kq�ֿ��S�A�����R����lW��P�,��P1��?r$/�����N�
��e��X���>8r:��T�έ!��̽~3���k�F��m �i�>��37_:lB� �Р�"�
��R��U�}��g:c8���j�l�P��j�v�p�@��/:}���P����6�k@�N7�#���k-F�̺Q;b��4�8?HKR%�:�(�J�'�~�O�c9Ew'�%ө�u2�
�JS:%X�.RQ��zz�F�(4t/U�oÿxsҵ<m�|��0+A<�3�WE�A+!�bi@���˗y��������G�7%��R\w��]�3���ÃG�D���ɘW�������Q}���n�J��wB������Ӫ{��A^��ԡ7HF�{M���$�}f��FJ�i[�~㱄�4gI";M `I��8$����F^�ǜ{|t�|_�fJ �6��Մ\+�V���Nz!ԱA�^�8�]V<��]�:K�mP��9�GB�Ƃ�H�֍�����98�C{�$S��,e��G�S��)�TQ��$�L��l�确.�J��u�>�I?l�GH�CX��<�2��%������?(�xn������!���[����'�A���A�u���ce �y%�k�����fO�`�SAͫnWҋ{�Ae��P��;R��"�0��R��S5��I=*C>)���h+)Xt�q������\��or�8����滪��ÏٻU��P��+$���t_�3y��;�j��/&�II�����jՑM;o!�y=�EL��>j@���jg�=�a�&��_a"\C;h_��*l/�!�P�Q:DE�2�EIڛx軷�Y*��0��'$��-��^�̟LM�[&�1�P�2�9r�{����f�7òp}�0_��xN�r'��!SoQ!�.`��}�g��A�}	���߾r�q�`L�[$�^�b��ޔ���[?c̮G
�'�0�ϸK�:i�13����!)�����t(�V(m�j��jX�N{4%�)2-Թz�ȷ|���B'�S��TfL�-5E�r���!?L)
�'�S�u�X�_QJ+�-��a���Ț�D'56��9�E�+�U�W\��2�q�����Q���Ͷ�1�u��J���I�D�=�0��}�A�z�k��՚_�&��'����U�[���!	a�
���iL����C�D/v��s~��h9�T��Yڷ�&z��
� /:M`og29�'�y��k�Et���Y|��	h<춁���m��E�K�פ_U7K�C�٬�ߚYd"�Sq�k ��R{oL���w�m4�~}�Y�JS_K����࿘����j ��k�]H��ᕝG�d7��'���!O�\N(Q�����d��	��WG�I��rK�7s��xt�����l�eg��ܲ�5}���������C��&��ݤu��|�ݻK͗��4������\Q��W#T��
������� 23�h!N?��F���o{�|����(dZ?�-�n_���x�hJ�O<�n�P�Xe�m�|����F����ڸЭ�?�^���{�l{��8��U���d�\��OXm�Im��H ݳ#��IޜW(O?T�#��#��p��{y!�q�c�e[rL6������*�	PԲ^a�����Ԭ�ʢ7àgUEô����� W8R�7��q֬o덹2���9���0)I;ВS��~�쵺���U���/v��8��	os�M�C��f��J४W<�F��.��7�:u��IL���.�=`�`e73֎��gIg�uU��N�o�&��*�f)f�/p)�������}�s�b�F�zB�q�.�������U�@��}���:@1�I׌� �ඨ�n 9��3���͹GZ�%���~��k�K	.���jX_�I�۽~�y;��ψSA�ޯ�1�sޡ����s��l���~u�V����j4$G|�p���/�հ��Y�&Q#��7��3�6HJlW��s�� ����%��)�UI���BU%��8jN)<�9:)
 ���Zp��I��w���.�V=�N�s������=G�p2�U��w��(R�j�(�j�j;�_�iϘ_�^7-�7H�'/LzMM)�a=5j�� ��A;��ɠ�FM��3.gvL}܀"�<����GbTsm����:�`�{���oSR�LcW��ʘ�{c���u
�%չ'�1�;B�>F���z+�����\�%�-�w���dv_5�|}�Nu�'"�$��2�y��1�<���鞟47{���,P-c��v����������
�OX��Wd�m�C�'���;\�'�{ͼV>���Љ�����lmlz���ϲ.;>hΑDu�槖&U˛�k��˟Re%A1�h��{<w�.���[�ZD�������iw�uR@�PAg��|w���s�tW��L��'�o_���;<|M�It_C�p�\�r�'�m��}�z/�Q���X 2�8���s'���_PZ8C>+ȣ��C��9�D���O��;M1,j�`I}��Y y�����жù~�3$\f��՗x�5�*M٤�.]�1g���8˹p�e�yW����v��{'z���'&ռϝ���f!r��6[�Ҙ�u�)�ld}�[�&AnJy[��i����	GB\�CZ�΁ 6�@eQ�O�g���&g�Δ�8��B���P�{�v�#k�T�jb��}W��7�u���L��<E�fY�FP�u����"LO.e�¸b��/[�$O#������� ���Vs&a����ᱠ�-�4�f�O��N�M�5����ݐ�@�b��yC{o%z�'-���=H�a�������@�@K�-�4Y~ܴ��eHJ�H���C��8��H胱�ȉG(vj���v�{�M_�{*BL��Zrv�(}���ۥ��A��w���;�l5����Ԭ��0	��?g)R��k�9.R�=��j�UVs*'y+7X������\��^H����d0*��g@�Z�2���
%r����:G;	U=��
�;�uK�z��x�.
�������X����dd�O���<�*Rn�j�ẶW`���♆���eҳ�u�}�K}L�����C�?B���Q��
�w��a�A7�t���E�l����SF_B�݉v�l��j��blGx���~�k�zݨ�e���a���Wl]�Ϥ�j���h
�tS;�ko8�YXKI���	�C���F��}Ѽ«�{��Q�$c����y��e�N�!�_ҝ��F�$�[����0wf��z'ʒb���Nȵ%W#�V~F���A�P�Jj�ƒ�X�Ps��Ԩ��9i@�["Ԍ4]�@��g�M1wO�%��#�i�H��/\<�Hwv�E����C�	e��.���&�Q�
���j�6G�E>��g�_Е� ��4�"���vҋ5.�O�<�.vr�p�	 ��S[��Ӥ�OD;�yP�[/��,�xQ�2$����{���_���Re��@xFr���;B��W5x���������3pHN-u������UTgZ��V}U�*ŕ;J��VZ�$%U���b�[ܔ�]"���uI��'�	Z�j�U��OX���!�|.�麤E޿=A���^�s<R����ʃ2I�E
��*q�����r�w3m�w,�W��L��6�����l�Z��'��\��V�'� 7��A<،COc}~ǡ��hK�񔂛L���MU��{��w���#�T#�߲E��V^���ӢV�h��R�\�3;�:$���N�
�;%���ᰕM�O��V���	��&tw{"*��yK��lP@�)��p,��ЍU9�W��P4K����珨���wÍP��1'Ko/d��'B�P�\|D�Yw.$PO�YR
v�K���[:�7�]�m78��nS�]�R���A6�=�+S�Um���F��~��� ��:.Kė
�38���l^��o�b&:�VZ�_�=�^'Ȓ��^q8낎c�Z�k>������zuN|:�Q o�?l�i/8�������s�a��fȷӦ�D�+{�23�9���4�7�e��פC��٩A;�k�2�pؖ����}�.�����cT����Ν�r��;�@�p
���TXq%! ᗘ���sd��Eò6+hE�+2a�鬚�?8q,�䒢�VΦ"��Ǣ��LO����=+��au�{�Xȅb�t���.��3���D2��W��]��[�=m�|(>9��&A^��K3���_��h�z�0vC8�E��T&��G��c^�������w���O}u���x�6����f�^Yv~F�t�EƧ	%�f�6Z�e��
�E�ţ&�G��~�RSWz���@�K(�k� \��z\h�tz�@�V���r|��1��׈M.<���-�.����9�9i�����\-�H��a�b���OBM��`V 	Й�F�X��&��n*	W�/�^zOI��Kq47���&�#��j�}�C��{A�O�6���`�<�][�?��f��}Y��k?xfu>��b�,K96��>8'1�W��h�����;H�B`~�؀�neǸ�R��j���X�S$���m����.ʉf8���<^C�o��^4��������>4t\��H�gs.\�1�r�J�Lz���X��.�l�Ƨ��-��]��)@�C�����}�y=���6�%y?��ve�X5�n��P:	M��ڝ�j�b���%�-����C �ƴ}8�x�f�oP����D$�ü�����JA�t`���Z�ij(�������D��}�cE���-I�v`r���Gi�z,|��Ez�Ga0���?�Tj	?������b�Չ�O���7ٹv�@yxA� ���{�C�������<KUZ�	9O�X��x�3�+=w�2�'�U�W�rœ}�>�� ��:�r~|�{q�I:�c�ϩ�j��p7���P��;���`W��j�i��]������XR萱ǋT�k���h�f��ό	eIϸ��`z[n.�r�3�'�����jY%BESҧ��E8ZDMoE�Ĺt~4x���~���+F���{�ܣsϳ��>����%�>l��WF�	6�W�`�z�P��B�l-�~�S�mYDقW���	e$�֓Eg\�C$Ө�p�DkMS���y��'�T�I����%�G��c�nލ<[��b��w�O� ����@(����Bх��ql����%<ƛ&L�Nc%VH�C|1�0�E]��MEc!�h8ɼ��T}9�;Gq���u�q7��(@�p�6�%�����}I���bL����~�ݕ�D�i��%�tѕ�*�T����83���­��֣R-�����"�߭���{`G���'��j)K_1�mk��Ej���ӢY�n�-��*Q�2	��X�s��e� �m7h��.y6	�����>hJqJd��i@�C��[JoSr.{1�k(�K�S�E8w��iw~9d�6Kp�m��Ih�N��e�z!����p��\�J����_������*M��zG�Je!�P�<�7 2d��%{�˄~W�=f%$�@������w7�B����V ���ގ<����ǝ�7G� �a,�\�Y ����lp|��R�\�R�2}X݄�̕��v��0/���n�K/%�����㷆��%���o$Cէ���Ff��'h�Y��dӉÍ�,v�#Eh�ǾƝ	ܠj��(~�bf��BP�1��s��Ѐ���(;2;1�,��\v��~i�цQ�C�hZi��GəZ-(X�d����.�OԀJo��K�"Mn�����S
���%��B�;
v����g5z�WL|�$Q#bψ�j@�hM�^do6k�d�M�t���R���.ܮ®JO�K*�e�lE
��^1�!�5«�tdn�R"nŀ��c����^~1�>�Rz�E�	��g�C�Q�q%v��tP���p���F1�;n(u���:�ib,#Q4�	:j���^��t����% �T,�`7����"�vm�j�y�^��Ģ�P;ݣ���3mΥ��q����*n�}����H�Տ<6�:~�Q�HpA�VK���j�蝏�&j�x�k�$�����f}z_E;�X�s#����<F�6Sy���4�c�C��h�T[�;�Q��~\�A�'PM��״�0��4(>��������?	��?��/{��s;Y$ �#8�{��#F)HN��+[#��צ4��������Y9��03f�&�?K���0��XF)]-H���bx�<7�/���Ǜ��Zɥ�%q"|�z\�:�ڝMD㕱���-'�H�L4�`>���\�(Q�� ���n�"�Eʌx�,��I.�*��C�eU�GQ����G�g8dM���!*ū%�0�I��xBz����h�n5zGVo7��m����d�v�u���c ��ȣ�$ʴ����ڧ��O�c�=�B�������TɃ��H���"��G޸}[��ߌ5�����o1\�j�=eUE	6����Mn�L�R�>��4��`�N��cj⮉��[e�L��P��dܜ�O�R�Q��3�܅K�PS�����w�B�,�X���۱����e�;�i����a�c������$R^�U&�v�)
`D�Y���t���%ѱ�]3��7R96�}�N��ŏrI�0nj�WjX�Y��ɋ�DU��+�$$����Y�<�r�*�"��-�	h=�8O[$J'5Lc��Ʊ��D|�����S�Lo��(Ď��=$�$v�W�T�����7�{�iz'��JS�ו���s��^�q���u�h����Z�=/�;@�vt��a�%�=._X!�3��´��I�T�#��m�d���Ԛ?o�ٖ�=R�,�����v�FUӒ�E�L���{S���g���N4A]GMv$�l�,�]��a�C������'�2PA���Q��џ��m�a���U�rCN��ZR4��s�D��n�E���������W1�����9yz=#���B#n7TV�-�C�K����@�U�����8�*�G��KOFKMWdYk��
�]�C��o��󽰽/@�,CO�]S�T
<�@A��@�,���(�fF?){{Ev�|�_�u	`kC�c7!���J���q[���ǲT��*A
�G�cD���)>lg&�F����Hj�  �'�'�O�����G���~���gʤlf�T�&p݌)��D�Fҷ�Fӿʟ%�h���R��l����i��e���x�`�ю�lET���mO�C�Hҗ�N[\�qЉB���9y(�*)5�ao��'Kn�T�{�<�īՕPYQl�.d>��a��&�ӔN��([\��>��ҥ��D�b�7��!��]1���~0��!�>Dd"ku�O��p��=�u����6KHS8���|�Cd_-C�i�mu;�f��ۭ$�W�d�*�tg��zY�7X�0�Ů���%���&f�|y�004��َ��lj���r����}�)~��L�!�	�`s9�:�i�n�To����5(zF�i���HQb`ˉ�g�tv_�`���VL� ��Tp�NleM�jV����n��?c���$�X���S��\�[t����n"���[����j�nD���H����/��U�D_��s݋H�`�Q�u�\rXg9,_S�N�9`�\Z�+�-�u#ҹ�fZ�����(��}�&��\�!��ߒe�+�4����mE D�<��&��sRO�0%웻B��#����Q'%��AZ|_ǫ;�`���뱏�' *���"Q�"q���3�=N-!%s�lD������?�-�MS$n�4�1nfxIt4ߧ*�X��<�%�w6<ݿo��X�a��*��m1�5ܑ�!����G3l������3��ҁd W�����I*3�#��l˟-j�;��T�C��@��T:h6��Z9�:;zt���d,v%�'N_�6v}X����U�F�K�U��g5'!�����IT ���p����؆�D����7���ų��#�8�\ck? ���+2_,� 0c�г
�@�\ez�����!�I~�>ڎW	@�69�:C�����s�yq����}n�Od��%6����$��T�a�c�f�Q>^ތ"���p>Ս8���J�)?������=6IN[�{���#1�H0�Y��~7�H2/�M'&`���<b`1�y��.���V�`��/9�T5'���(j7bY�'���؏����E;�@R��Ӏ\��a��0�%�֜�*�>ŭ�%�*���1���"�#��'W���ǚ�����u�~���V���̡P���r��݊��|�c/�M-����]9��$� ��[<�Y����o�}��lQ�ʞ�2+�0F�/�$쑲�N{b���3\�ͪI
L�jw�#7����{ ��2�����J?��ƽ~(㺙2�X\.��)��"�"I���DH@H=�<�n���]<-=9����g<�uR[^�X��X��\~�泡�Re6��w�e�P�z�a��h7�C���+���W^���O�>���&��!�!l�lN����ԕ-�<t�����o=3�D�K�R��O,��!��m�EC8�չ��7��/����yW N�J��?�,�O��;��}@ڮ��T�tj7�㬑�ɒ���٭��]��O<l�k�`���2��i��9�����̚r���<J��{��Q�ÙbvS%�����p�\�xAXj���V_Hnpc�ˌ$�isn�l�D3��ЀS(/�?`�ߒ^�G�
��엍�I^���̕t
CC��J��|l� % X9�x�؃�X':,�� �� �e���}M��w|ﲪ��7�xy!��')D�3�}�6>�#����x�No����dV����.�S�k&Ң<J�����C��N��� �ͫ(w!�=��G
2��^^��`�h��[��Y�����[
���Z}'�>�8��I�#䘷z�༈4?�ƞ�ĴQV'� sO쳹!_օp��S+M!wG9��|'�fʨ=��Hװ�HL&�wW�6�5�%������I�"V@���2�>#?��y��9��G9��ސ��4Ɏ��]re��ƥ8��cK�����(�����-e����߆I���h��ԫ�y��"���Ĝ�V��M�� �@8���l7��j쥫B�o�;�P�(ܓ͛��I�A��lm�@@�v�}I?��T$eR�2�q�ׇ�V�z7������D���Zٽ��i}�ς��6j| ��d.�.��+���i���G��f��Z�h¾�#���|�E�Gz�ǌk��ٳMi��?�����o�?�SMo������f&���eD�8r�lw<�]�S�~�<�3�G��d�.E�Z~�!���q۩�~��u[����|_��+NQ�.):��`[���e�h��"_GlbQnt
x�+���㧦T<Fs~ ^��k�P�:�iS��{�FׁZ��˚6�?�������O<�4!FP���YMx(�ܞ\޶�eUY��gD����R�p�j���ǍI��lsNlfox�{���H���]�%�7�J���ay���n�$�/��r��Ō:3�k~"����d�a|C�\=w,��Z~
��>\fB���BE�'��������c$R�9b_�5������� ��u��''�tQs,{�V� �xYI?
�k�Q�i8���� �,��By�!�D\3S�>(ѱ%g)�`�b�C��{}b@}�������䥨�H=X@?[\e5�8�^!��KY����cʀ�xrb?�_�&[~PtZ_`K����e��1��ZK�ò�nŚ����2��<���ry�s�@��ӏd�.�>�E�����YE�Nߙ�q�<jZP1 ��D�������?�:����-ј��c�q|k���E�v�O�=4�^kB��3H�lT�+ꏯ�c5=���Ə�;��{g�׽f�a��N�	v�C�<sk���d{	o ��~?˴�s��������8�v-���Vv�q W��7�*f��e�"C.gq�2�K��%���?�*�"�e2L��7�Q@y�9A���Y���9N9X���E�=�]kJ�U던����\�yÜ����m~�6����	4d��J0�I���2&"%�ԛ�A��+8������E��K��`��B��}���'?�0J��ڲm�,d��i'u��#��5��`�g(�Bt���N���I~+�
#��;��iI��tr;��
��z��厼�e�'��w���Xwi^��B9�����"�j�E��xpG�r,piN��S��v���㍠l�l翯{н�3�$P8����YR]~��ӟS��»���_w�n�PJ��GP�#���x|�+�>���+i63&4`�����L�����?kh�p���U/�^�[YA"�k�鄓˩mՂ<��L��?'����F'5�8_�= )I��$�PZ�|E/��\��$G ��#� _�!�a���?�5i����{֠�N��ǉM1�6�{��S9_|��H��x���mOM���̧�*�>���=��*���q]v��P+��tE^,�nO��.���Z�
�5�*ɬ�E�|�ZI��#*	tp1���w�����\ZY������P�-�/�V>|')���K[�n��;��QY��繡�|��{՘<mq�\�U@{��$N��ꗭ.D�>�b��(�_tr��p��Ŭ���r�n#���4.<_%-p�5��=�<>lx�9Q&���d�i_"@��[v~���'�Pd��g��L �ea�(Y�*s�~���/ebB�J��1P�ήJ������o׫y�1�7�l@hlP�G�`�ԁ�@Z��°U[%�����w��� }����ԑ���&�>��6f �$�4n�T#D��\d�����;��&/0vzD��z  M����&_5��q�߱����Q-v>zl3���BrJ*�9�ġ��3�'7�W�w�Ӿ���ħ�qx�֙�}V�TQ'�DV�XA�K�p����)M��3�+M�0��\�o����z�������K��
QS�+:�hs�1��R�f��hx��������Y/	 XNJъ�}��g =G%��K�,��u���5n���K�`��L	��e"'����u @K��U�Qݲ�'��a�F�Q?�m�ֳf��D�(��s�%��bP	l����vX[�����3�@,���_?��*�"7j�F���������BR55/ %g]�  % �>�Kq��f/�G'ʛp�)�pRl��B#�S��ɒ�֒�-"���O�mV��g�� (=u��)֮��`��i�8{�ㅷ^x����Dn"3dan+j`��ٲ*�r0�Z��~���<`��瞶��+s��U��hi�n�H�'�k+s���)��T�V�GN�p��H���)wI�|���l)�!H"r�ڍ�:����n�q� 3�:�C.���w>qw�!Z ����
���������J�����<�W��㶉����ʴQA�o��3e-A���r\�X���YY]?�����������ͩ����I0�A]��w�m4q[��44G�0[��bZ�O��n�"����%i;��mb#*G~�@��p�C��>U��M�vX�g�Љh7���1q��n�k������'�8[z�6�8��	�.z�k�kiTz�M�>*��|��;��I����d�'i~;���Q�N���/��\غ�����Uc��n���K�s�uق��WD՝ �lļ��·���Y˸��w��<�?�!�D��E�dx͕�LUO�礡�1�6oŬS0�aW밯�5֔X��8m���WBUu<<�$-����<�	d7	��5���7�j��Pq����0��`� ��=��5F��|�����9Ɨ�/o�/�`�1�XJ��3�n�-ţo�m=R_�pR�ʖP��<�b���;U'b#�:@����b�N&��9�w�7���V3�|���j��'S��� {W�:-*$@��5���i\�1�f�+��ֵ KSHR���ŖRlI��:�p�(�ψ�|6�(C{���I�.\��rVl���>��{�s5�Qq�H�A���[�Rۅ^6��0v��>�"���R4����Y��f�$�R�sk��p�{˙�$�w�2IS��Wn�~R���a���Ǳ��S���Vl�/$'iC�5Q��xq,Zf�(=�}���� ��yD�Ǥ�;P��o��\1�H�3N�����GE�����P:���Ε��J��\P�csG}չ��$j�ܓ�>%ZD�Ѧ��=�6H�����k��X~�����HԟHͅ�Q]TEƜۤ����G�v]�q�#�����XIx:"�A<8)��ʻ��΃�N H�4���4�?/��_�f�ίH�����}]��Ĺ�B��,��+�l~<�n]
\��Z�_���0*7��$e*��%BFP���^�n_�U�7��hb��	�J����K���jF��v!��W����(�D���
��>>��jPV}�ԯ`�(����yrV��8��) '�)	��u*e�G�� f��-��Nx͠�괇"�Q�Fql�����51S�������~�W���2�n$�U��{�^�PP���?�;ns��=�~_��*�{1��yJ�����D+gQ_���������}k�۬5������6�1��ؾ�CP���?�8��4��$�����V��
�o�6$%�&eT���fvz�|h�ϐ���|9b͏�&�l���#��H�����4�o��\m�~
��FNv)�a�b䜗��E���҄A�x�Uc�f3�z���{�Q-	�z�����`��lv�׏A����د������V��N���C@i�w`�����#�� ӂʋrˣ4c���?G��E+�o(T��P�*�tP����e��j$2��	sH�$�w_��˓f����t1>/Ք��������;�F>�Q���8�)�{�i`�x�3^��ĳ	
�h��P��K@����KF ڸ�m[]טS��Jl9���ha�g�n9��29'�7Jn�yõ�qƲ��P���#�O��Z�k~In����0k<�(h�����ޕ�h^s�G�\��v�NDRbo�kw�0��H�e*J����pTQl0��x�Ⱦ�t7WU�=��xR�:e��kP���4�3Q�U�EZuD��p�߱ �t)��)B)zZ��e��uh��AZ�y��1u��V�w��ŮO�����:�<��ekT똒յj�f�Q~����]���W������ā��}�y�H�6*�r��,��Y��'N�M���[�H���y�,\O{�U�i��|�;���f�0r�H�2Zw��$��X��kѪbbd� �B=�����+�"��'0�]mf���H�Z���u��
�$�<�őԨ�Zi�nc���S]-d�1)�R�K��)D.��Lu<�%��Q6��on�~�7q�&;,ಈ�诖W~�������J��9���*@��ڜ�`�y��P	�#E��Xm�<qB11W���[��olǢ�CQ�	���j���p� �������;�?ΰKwؐk�����Y<ҏ�GI�,�ף��]m����D��\s���c��[�'K�� ;���]Y�OF��k3��Z���|cUI�W_I�65�=A-��jVZ��j�w�A��c��=��e^��Ք����XF/Pf+�'��ck,1���M�(v9S�j,9�[�7���	+ 8��8�l�7�@@���U|��/ʡ?V�h./�W���j�E���cC��]�i.J�/�ҍ$�F.��Z9��矮��[<���"_+j���見8h��;��kWk���қ:�2�<�K�#���z�sr|��M�op���������g��*aҧ}֮���ũX�+�4��hg)�s}�|�������Q%�߮x������y�u̙�G�L;�($��M7�s[��M_4��j�����7���E.�,(4���v��� �M<+	\}�ӣ�����h�m��!2;�h�z���)���)n������Lh�ܾT=r�}&�7B�]��j�t�*�����*0�?��l�(6P�;�h'�Ơn�͡�=n�P>�-��c���VFҫ� ���U4�'��1΅�߳�(8iO'��e:Us:{�K�۞�a0�RRn���6y����ߛ-4��o9:!(cs��������QǌC�J7]0� ��U�Qi֢���H+2�ї?�:ߏ�+ZEۆ�u�t�+sbMD^���ly�[�� ɵ�K .�58�an���!HY<&���jIx�U�JW1��Ъ��~��J눽��U����#����B#:\�l�ڿ:�֎_��3�ZpE_�`D��'6g��c��S�]��yy��3 
.��áͬC@T[,Wү��Z�����~>�xfgI��� �FU� q�Fzi_ �^�$@�C2�N�S��(���D4�w���B㻟&VT=&���|�yp�A�ɼi�AR�'q�^�@˅���a_�zl&��T�{�3=�!�=����n�$���^7?ʿ�z���9��泤����6/+;���>�?���;��=qmm�I�m����3:8�:��o�3k0�
�&��d�kEm6����;}��s��_#��Z.^�J?7o8�~��I6�X�ve��X���|�x�����r&�a0*&\�O�z�4�����|}�M���Rۜ��f��JE�P��\\Ι�	�c���������mC�G��h%~mjl�PRX�L&�������1; ���$�De0���E�S��^OG�Xܔg����V�CQ)���ə�¨���5��ezЌ8H��n
�LU��S?�%�7�p�����	��>�6bh9�`'�1�7WuU%p����_r��?���	ϻ��5��>�!���l�1���u�=E*�갋>�.�����
��|VE"U��F��z`Gn����d��s��y�f�A���?x*��:���ݻ�p4�������������>��#q�	w|3D1� �Jk�����O*Ρ�t�j���s�m1|��JDs�8\�nc
��7Q�9�|,�+���eNP�^�,�Y�ռ	=Y��|��פjDW�"��c!���]��ui.b��;?c�x"6+�u��q`�P�"7E��8%�YP���Ѓ���B���T���3,3�J�3��]vf(lk�7A,&d����q�7DP�j��j�0�l�^�]�`�Ś�`��w�ƿ�k���<Ri1}UB���>�?���b'!7����/�`"pW�����&4�tՔ� ǅ[	�o�ʖM�"w��j���1�\�2�"�A�kȅT��G-����MK3�Iμ%D�W�U�Q��}��9 B�-�ΓS��tꞛ��^y�ރ�����M��?����:���A�p�LG���d����ľ��ӂ����`�B��a,��Q��u�FK���1�����4I-�]�F��t���pI��+�����ؕ��%�/I��l��� ��5!���UbcsQ�x�eow�Z��B-:-�B�A*/k��hE�Ьa�eU1�q��Fіv75mv��MT�t!�t�crz�tc����)C������m���mU�k�y	�+n��s\�Py�_7�L���s`���muF�\5��2��.ؗ'��:[!��7��m�����A�l�чKj]s�m���L�ό�Ȃs[��<��$�0�ج������@k �� �O(�#!��ts�3~x����r{��؈�.���%ܘi�k����\yt�G~ef��;���Rԋu��O�Gz���9�����N[��$e����3��-�Rp��S��2�P�5^�m�/6i�Ͷ�`�IE�he��)����̰���=M}���XS�b�F�����%�ܬ�\`�6��R���������O�ե����ϡ!��{�Xq�ʧ�0Dv�l�紳<��x�9����"���gW�m
3�u���c�-�#��c�wRSmR�Oq���ڧ�J>\�F	�}�,��b�^|?~P͈WWj+����ǟm�`�,a@O�!����\�NG�����1MϨ*�lwJȐ��a,U©��R���'�\B��2�}����O��(�>���>0��1�!����w�O�	E����_ �[\ZΊţr�
�!��ÁX�[�1AQ��=�����(w;��$�������-&���v������6�y�V�o�&��<��ܰ˘zT�+ �a�(��Du���Fx7��o�q�_T���r{��~���z b��l���츭��V� b��>��G:�� ;'���@�1�h�UǄP�����Lb�y1
3�-�4�����0C�C�=Mʲ��j�/���l�m�/��-LI���M 9�d�7�4͓#��L�&��|��S4��0[N�ր��H��УKԏ����EP��[]�7�(�Wy��S-�;���)��E2����F3N�ժ�>O6���[B����8�;ϳg�%®T,k�av��"]�$a����1%����B��np��n�ؽ=浊��1&t�
�	5גZ2ڑ�xvT��8zd$=����{Ĕ4A����dk���m�&`�aXxp&-�	�뀂ٰ)Wj!(X�\+)�$e����ONy�(��:$��n����4Im~���c7FbO��󇳌�L�n��Ԃ~�3���{�F�� V�Gr[��C��"[%��{�T�^\3uj�G�K�Nצ<�s���޼
�
��!�GN$�Po�p1Tf
kV�����uH��z�Fυ�kHU'���E;�'��X�|�U���Fڒ�rG���p�gEn��8��:���
� �Zđ7�]��!VR��A��P��cx�r� ռ��T������z��~�[l��(����*�
��{�!NҲc�OhQK8���]�X>�b�� [9�I�[��?\7��`�?��kD����� �Dpd���D�����Q�6v�d���1P��
�rтq�U�j���bRy�7T���_�wɊN��$�|�˜Dq�Ip�R����Q?A�5*u�
�A����p����m����W؋���Jf��ߐ�A�+��i�/Ρ+ ������������:1��Ol�d-���������N�����)of��􏘆]=���K�"�Ϝ�f����T]n�Ǘ/m���]�&���>+3��,x!^6��냹6����� �r79��!���j�&i�B�pD��W��Z�$�]����h&
��F5�V�6�e|�R����1O�FO��Zɧ��ۤ117f���5�}?���s�	����p���%��+ �;�ϝ$K���̓Q�Pw�"����7��V4~��٠����vqݹ�^J���.�=}�
�`��u�Ñ_��� �`
UU�0MM�a���@��@�j`G���5-y�}��m�>'˕�Q赲+7!;�՟/�e�l��n�K5'f5;��2�N�ѡ��)���@��1��(�,���?$ӧ�W��ɍ�ɍ��G�`?8����+%|���&�G��I�J��zUd-X�L�c�La��O�!���\-�m>T�[�+�?�=��蛱�ݶ�9�j�����m�庑(�;}�,!�rr�t�( ��~Tnz���~�`!	��ar$�]���RJ���R �S���s7��ٹ'��#)�#��z�ח���NlY�P�H�����z�4�f�/[�ʔ�IE�gF3�	�7<8O4z��"��PG��t�Hfm�G*;������b>�6e
`9���|�1	�Qڮ����mF��� ��}_�$���}X���
y���՛�FO�Na����.��pLL�bp�����W����9����`쇨fM� x6���ZEEX�nh�S�{��I+.~Fȍ7.�W��*�=��y)V��
�	,|�>`J.}�Z�3�Y��,�V%Ri�`Щ����k|���b�y���r�V4��74"���fxg��aF^x8�n�K�=�jo�B�<#����/J�A��c���`�m��K>����A�ғ�X�i�C��т��^�ڑ�*h^U����w��������<���Q5ֶY>z����\���s�#������^]�6Z��CoX�]�\w�`X�ԟ01j.�S8E@Y��յ,����F Y��J�E�e�w�5�)\�ٔ�܈Lk�vA��N�Ћ�����3qL�8��(��҆ǁѰ ��FGG�vv�|����񺌆'�Fpx3��6`�-'y���^�_'مk��􏏣'up*F�rA�}��ߍ����eS�Tn�c=�M�a����4є�+��]�����O2	ܮ��cTQ]��-�*K���Ov�s��|��aه<����.q�hJ_�v9��̊��QS�eA����yQw����߾T��w�U'��u�FC�']����q���v1H�V���;��3%;����t�4�HR�n荓f�� иeZ6]J5�eŇM�7\@��M��q��V.��Fp}ӓ|��-�ʢ��B*!��Hz�i�Lƍ�����u3�
a����rJ�J�z ��K�n��uE!��"y��K3��s��.��$Zitt�2�挚u�M	�d��̸~C��QV&޽E��Wć�-��|�l����i���� �^8�3���mBg���<Azg>va9j�����=��N7��<m~DϢB	W�gv|q����Lb��i��q������8�sᵇ�9�+���%��j�Nn캆a�IS�OY�5 ��-"r�(9���<wl�J���yRe�M$*GC����N�o3Z0n�7�О�\2T"�(r L튝r���0ެ6��l����!�
�4z�(���[������Q����
����'�\��$d���:Ͷh #�TL�JYd�hO���v�����M�����^k�ƴ_����h�Ɏ!��U�ݖ�F���/��ߛ�Q�u@�6��]�S^��Ž��.f Ł;�g��_�r!��=��:��1�F�:}S3-l6<Ŕ�u�1s4�>��9�l�!v0�ޱ�4��V�H���[OPz�6 dZ�,�x6��ga�'f� �w���� �]���o�&!����*#�:�\1��D���W�n�5HS��8���O�.mjë�;�I����.w}ƩGf����֤ �h/,���cB����C[R�#e��!3��U��E'KJ��*KU6�
��m'_~F�I��D����یGS��y�J{E��}R�nz��%�	H|���xЦ��A�=a��e"j���U�{䒢��F�I�G��끷a��YN�F�E�5p��1�5�!�*��I��q���t��*�B�I]��m["	��2c��d�
���$wF�]��ש綐S��{g=K�N�x�7�v[�f��3; ���XU�����_�����VA��/�4��D�[���K��ː��	�����ļ|
YL�Yq?�-`��L%�}�s�f�%8����*�EX*9E� �E�x��Q����S��c��&Lz)���N�I�~��M�ڬQ�H��5��	_�$��-�T��]���)�ݯq��{F$6T�Q!�MmT�����e;��{j���݃���鹶�X2Ԣ#�#w��_���^��i9x�PW����Z1�LK&��쑚��h�YO؎jVHf�L�`*|h���� � �f�xf(,��dֽ^�[&���ק7���o�9-��0"h:������R!)��&�-�:��E�;���2VTi�j���o\00Z�G�Z m�C�?�K�\xF@���0�7%aD�ȹ�`[(��R|����jB6,���P���6N����B�?����
a�F�g�ԪϽm>�\~o��z������e8.���˻y�G�u1��Te�
�2�����K�(���[�"�~/�P� S`��)S��W�[�`�C���0ث�S�o#N���^U�4"��X�,�
��g:�#	��r����n�F+@p#%Ԍ��Q�#n���t6a*�J'�Wd6!��1ۤK�꫋����2�%�k�{��Y9��#o��<�z{��T]�;Ԓ��J�&P��e�NꁽK�X8ʂX+�]����Å����M�"�������Qs��wE����YD-A+K �VjJ/:�t��ga����W&܍b���@M-�#O�P�g�ʋ�)��i��;-�J��P>�!4a�ck��g
8��g�~��<g�e����5�{��d�4J8I��mK���-�Q�#����$�7m��� 0�Ҵ7r�6d�?0F�� �71V�V�h����FgtdTΕ���Ό�e�dv︎��j?������j�:�־�Y�����zJ8C��="�D	��}M�&ʼ�彼�"q��?�ۄ]�ڒv�ͺ�4.�c�V���Q���K �秃{���>����Ĺ����`i^��3��X�dY&�>�O,�1���v����>��������� :�<jA�!��:����I�[��V[��e��9y�`��<.�>)�5y7��7�bz��Y��͉����I�:�QA�pGD�S�뢡�E5T�J_+Pਮx�a��p�_➑����ޠI}�
9s>to��!	��J�0uyWš��c��!� �[�J��\p����@���XŬ%C�Q�c� ���rDO�E"�@�2���x���K��/�p��H�� �V�
�g4&�Td��>җ���C�y�Vhhl�?�t�_�>�ę�;����J1 ���.������$�}3��)��t���˛�vkc�?D`*������~�=� 3SA��x/9���
+!�U3J��ku&��"����q�z���K�W��+����u�M�z56e3�C�D;�5��ͩ�6�����˕]%�Q�
q|�s��ߺj��aԲ�lK�Z��?ق��ò�nۧ� O�r�t�Ӽks�&3,I�0^� i �0���0�т޾Ar�N���1.2Ń��*6"E��O�kQ�%���^� >�r�R�XM&��M�QpJF�&�~�{	ce �[W�`�
~�0_�ad��zlpp����!g4�Ӊ���03=�����v����Mgˁ0��5 ��(3�mf�� �R�0�X�>�JdO��ðKR�dΞ:����hJl����^(���]GR�D?FM�ZWi���|韮��7=�j()����q{�s�h���\ꙕ㠸�R��.{b��m��c��g�mq����t���W5:�]lG(��«�V�i
ϵ@����<�.�Ʒ��K]������.GaҼ�f��h��d��v���~a��kn��$��x�G�gC�3I;��R��r2�쥬K�&�������C2���0��9Q�$ˌ~09���Q�"v/ş�nF
R�1ck0�����^�0o�ӳ�:e^�E��3��0.%YP��쥩��/�HD��rw鉭쭕A�b,��6C0+�	Z�c:��ۺ�L�u�5��tӳƣ�PlfL50NQJ�Yv%QF�w���*�N4zz�߄��,�I��[�25�U�.�ȗp����M�=� H|��x�<�j6z/X��:��X���e��lK1�c	��'�Y@BܦXDKü��|���-tr�.����ĺ}����Cp��
�V5�ą��x#D5���IHyo��@�g-
n+)�ҷP�T�&p(��܈L���WU��ւT.WsD}�U5��&s�Z}ktB0����"y��������I �ҩܘ�w@�9�1��N��櫇f
S�i�	�����f�� ��}!�6J����'� @��І��nU����	��8s��]UB����ʲ��n��v"�Ux��p�s�A4���ȿ=��	� ���53�
�k�Ba���B˟�o	��,�Ô*��tS������33l��N��5�q��Ԏ؍k�X�Q��������u#���N�L��j#eX"�&prN��NH�ŝƠٖ��E���7& ;\���et��v�r�i��O�ͳ5��@ȱ��hsỬC"�(
�[^����C0j��~��f�$�nʎ�=���Y���Nqk�pA��nP�_"���ť_��P��L�J��":a=�Q����;Y�&��3'�3����>�s'�ZA��p�-E�ճVJt��|P�ܥj���M�_�x�e��,<`��V�?V��,cSwX_��yS;4&�])"�	�)�c���W�Q� &��>K>	g?٣��8�>�v�"pޠ\�&k֩|�00H��<5z�
;SV���֪���{ȅAED�=W+��ֆV�Rd��C	W��v�q��Ch�+��3�<�(��J�3� 1�(M[������z�Y
�d��">I�l���!�7�[�@��/е��ׁ~8�W��
�R���FI���j�>�щ6�� g�����7XS�K�q+�7*�"�Zv��7.�/��WV�-<�	�^�gf��(�F�0bhӟ�pmA���-��j�``��i0ް�aB�k�I��/ƅ�=VsB+�x��]��s�U;q��p�J����bA;S)��ٝ��q9Y��Z�y�������/��^P���FUۨ���(���C��w�Ѕ�`Z�}�_O�ޞds4l�?�:�˪J{$36Ι�!B��[�1�yC��D�@�#IC�ټ�v��X�R���e��i�����L�%��3k��F�Nt���Fdb�C�+a�"l�?�ׄX_z�rV;~�3�ea�#��{�Bg3�[j�`S��PS�6@1|&@=����h�s�w��@y�l-�v��/r�D��9#�[Ȟ��D� E�l��9�Ҡ���댟lѣw�أj�$���4pYh��P��5��|>�a:  e�(�?`����	ð�{��s7��l�Bᚧ���a��e����d�?i�"%����ѐ'�1����k���xg� >}���:��R�Y_vg�M\UbRY7�1�l?�`�^�'���5��C\S�=B��0�d�zhsRɉ���s�Ќ9Y��n�z���
���fd�Q���>��F��3t+��T��۴h�X���4��,B���Wۍ����髿Y#��&>� Y�8]r�	>Qd�-�s�c9� ���DE(@7�u�pэ����p��:/��ܓ�klѹt<�D�[7��K���<���TS|��E|���\��uϱ�
e�>*�pE󗷒u��c�C�k_"Lp@��_*��~��Zۦ�4-���t�ʦ?���6����gm��e�xu�N�8��pE�#�h3��G��_�+��NX��/3p�|,��.��C*��pT��r��>{�|�����k�����0��+L!��ɖ�'���f��[�6�N"�/�ڙ����N�
Ga���1�?�ƹ�_���԰����a���UI�kF�M�;��mWLz�-F��␷��sҠS�x��5y2����B���{ɱ�9����\!7�yx�O�q�����3�GSH]ja#�dv�K3��4|(\��ޱ|O��݅+:ܴ�%����3��l̞Q"̥[h^��Q}��a�
lj��{�Pl@7 ���XB�&�O��Z�C�r��������G��ЖV1^�UU���8C̚Q&׽��p�8K0����Q���H\�|C���LӮ��:��S�T��.U�ՙ��H��Xj�g�a)�@�����Ԟ�L��F|�M_v��o���w1X��3���j$�FP5p㍈��"@���!$�ݝ����� y���߫ �n�ɰ���`�-��l�%��9�Z{h�m]�$-S/,�Y�5�9&* 'A�8b0���ٿ龕����u��$^�@w0ķ��-Z>�ܱ���v��4j8"��'Sy��<�&�d݋�����S�IB �L��nC��3�N���2�:�uU55ج�!(I��]�@��:-�O����#�� ��B�d��M=N:�"����l�+0Z��r����&�.v��}�
�K�5���%P���b�b�ΗP�NW�8Cp]}r0����%��A��㼺%}��n"�v8$��X�ӭ��S���E���{/�Ư��/<��A��Pũ��pHԲ�'���L�����Q۝OWN�`���Fz�m���X��k�r�u|e�\CԈ��
[�� Ȧ-�K&���tY&�+#>dE1�z��s]ɣ���=�	�jtR��pe��S�hzm"rRշX�-����(eו��dD�����v'��o�=����8�c��u�:�d;�����W�l�"���df�{ޯ�X��H��] �rnd�����!^�h&��W�
�e/��ܗA�qrn��l����TU��A�N@�;�cn�N���~D�g�=r��k��(Sz]��+�����ز�Q�;��V���~�6��!{���!��w6TL�q8.'}m%�3����dcA��5([�	$�_�a)�]�~��Ĝ���A�ɜ�X`���gW<���nd$��Gt�E$rl�(�d��^�;�����#C?>l⤚9�}�ˈ���v����3��7 �L �C���Sm@.�v�v1���3G�X)Z۪J��&;w����#��A�w�?0V�%��͔اqi#�}7o̎~�o� �8S�"�	(yP(ߟ�߱��{��KqN�d�TP4���;�Ď��s�g*�.�4&�I��{�,o��_��:�N����;kJ4���T��3<�����)�lʲl'����ߤ�.Ĩ���v�a�)a�<�p�y=�'6�9�9�U�_]Z�2��
�_H%�-g(�G���)����e@��ݍ���U�[�1T���(C^J�$aV-[�:j}v8+.a3� q��JCN�_l��T}��L�>�XJ�>���V)f4f ��:�Υ&(bJ��xuMh�g���~��/���fT3��6�:�Zd��&�z�L���]0clX�)ً�V���������ݸRy�~ǘq���Qػ��Uv+CT�m�ͦ�,h��m���G�	�[����Fvʭ%�E_�%q���!������馢�y2�@�fZ�@��+p_��=#���'�k"���i��eZ��'��<-V5�\d\xC8l@מ�3��Sl�v>M"��.��rr�������@�LO#�}#�ʁ�w�%�o>O�hY�i #0��Cp1��
�P��P.l��7�W]d"ϐ5|1%�,ce�ZH���J����߳�E�>}�ӧ��x�l�T�t�qy�!ޞݖ��>W�x}P�'�Mm01n)zC=�b��ǧO誺�wW��Ԓ�q��e�H�wr�Ab����*8/����V� i�"����s�@�����8(X���~Ζ��d7�h(����̱ZU�.������4[!������'��ksǈ��8h����L�t6��M���#��
f������5�&,���B��u7��<x4�Me�&Q�f�1R@T�mI.�'^�(O�
���k�#]�	7�����8��]��hz�AyoSj슬rnT�D�hB5N7hD�&;�'i���aC���H��NU�_!8E�ԼZco�K*jk�q��*����&5�`6q�Is0oңXv�s�<�>��R��B5��a��M�i�����N�vh�~��*��ڪ\|�bl�BL58@4�'7O�l����_�㎦�護���I@.�� ���?��V����#�{A3&z�p�ԣ�����Z��c ϱ���I����NE�儖w3{ y��bq��T��|��E}:����X�mRH�P�J��:v��S�
��?�د+�x,�k;�DL���&ZO%�̾X{0�J�R
!�h�4����p$��Яξ��ӫ�Ȯ,�Hw�0�FzvpK���/I��:�#��Ϸ�E^�x�=w�E
�dL?,F�#�������h�*��$��ǀ R5�c������KQ��*=r"��f>��|>Ήg���8��FmJ�^���&�r*0��d�#֛l��pG�i�â��+_����!ۼ� :4Z�K�xs̛t	F08(Z����I��	�᳽�:&jFƪc(k�Izoj�	�_�Z_:��n� :B��l�e�;��r9Oׅ$p)B*�]��ߢ�x��y����[�]�E�Z�Mv�Z�B\�M�����U��������pSo~�U�w�v	�*�����S�證��9SS�d߫tLj����|&��5;�1p�JZ&?ʡ��T�z���9Ŧ�r�|6�hl��9t1mm�[�]��:Vw+�Gq>���q��8:����T'��(�m&�^H��M묅c���S�aH�$�+R����߭oJ2�ed$��y�ȃ(��C��W7C��TĉN�L�:o5��I����[��H�zyX2���$,{|W��O�?Okv��G�ҡĻbk{O�5T�KI��������s�v�tQ%Ť�2���roR4:�f�vY���Y�l0S�BMwn9��8~^O�|��:'��ǌ!� λ�5"]X�E�˴��-nP
9��6�Dw&�x�������7e>����pՇ�h�-0�-�Qu,��H���yX=؝_	�1��-2m�ʨ�հ�[Lј�
���/��1^�Ʉё���.@]ta�i��З����l���)��������@0}<����x���k��Oh�i�I&�V"a�š ��D3#��=���+(Xjڿ���V���m�)���Uc�Y�U���4~;�k/憹��q��� �%ר�X�TX��LڑW^����Y�Y<��F{8�O3l�)�D��H*�}�˙���E�ݒ����3 /��Jr��W�p������0}���Tw��bE:�cG���L�!�N!6�Dպ�\���o�1���S�ZH0ȃ�%��M7��R��g�JH�7/7T3U ���W�r������P�'?I��ɱ��e�$�U���c�R�_��j;h���h�(ڰ���o��=z�D9$�M�Ҹ�lƌE�Q��F7�3�Z��s������Aև����h.�P	:�&�Аߘ� ��!F^W��[B덦��Q�0��&������	�B�?i#�X�Q]"2=��
����1��xQu�<PxRF�_`�*j��(���B�;�D�n�h�;�P��o�C�
΄"��<���qL�
�Z ��?�>5�d1���_�%�#�ץ�s�1�t�h���wPp�^+�3g��ڨ�B�k��~�K~�k�8q�ǣS����`��P�X=[�uoa[��twX��Uy���\(9�E��衡x�Q��9�F���Ź��	��Xݑ����y��g�z
1��i���/_6��
	��#�!�y�W)��q��*�5�b���sΌQ/^�Yr�T��]
��r����چ��"C���������;R�%���5��놾M~���X*L�����<�vNyR��O;D~Ήk
X���'�VYb>��E h�n	<=$DVe��^�F�c`�ґt)�yH��D/k��{"��疩.�}��W���vz(L�EW��3��12w�8��8�!Ԁ]�7��/�C�5�~}�N$}������A8��܊[E�+�I7��B���of\'!G��\��R��6�|QF�H�5����=�#��R��?D*r��u����8�����G֭^��K3����8-��^Mq��}W@
q�vM�T�uQu��;k��Y��z�4��Q3J�*(�nMf��?=�U��N�r��pL��*M�h�Oa�ܷ�;�I��rB����X"�=Y���H?�N걉`�������	�O�B�w-�9@���f��z���/��e�7��5���V�Q��.��we�0����$<��j���JL{t�<F�,���~�@�ҷMk��=ό��D#	��їy��/EO�;�C���Ks����]�5��
�6���	����˲�?�a�IS�@��?�\�(���pKF�w�������}����\��~��S�L��T��j�g�RH�%��{[T��Fܶ�mޣ he�%�t�\��V�>�!ɤ�m���P��B���-��BXm!·�L�;���ě�@XM���n�[���Rk�s8����]����eF2m��T��j�q���V���U3���0�?40�KL�/�<�r��$�[��3(w��<��A�r�w�Eܻ>��o63��r5��&�v�����	_:ְ���[	p��A~�^��أڃ�k.�N�4�����U3=�� ���9�v#Z3^��?�M_��I�O�����JK�{u+c^����Myu�S�_��Ih��A]��)
�B�
��O}.�np0�8�I����P{�S�ȧ�K��0��� q*,��f�X�|/�>S�y�n��>�p)W�����?��q�D�Zv^��U�� ������j{b�" I�*$�ں���T8�N�[���a�\�3�e6�(�vx��p����6�A�.lxx7@�Cn�)G���F �U^1��`����!�v��x�l+2�f� ����;q�m�=-��!B+��6��.ۜ��o��\۽���0� ��������.v�a}��p�=�t�B?����6�<�[|���a��"D������J���㘪j�]m�{}�Zn��6:�p��l�X)�� \%���4���w��p���\�G��8���9G�	�[��K�̀��yJS-�<�������OdO�H��賂�rO���Ch=:{v�|�ZAg�=�S6��:��x���w
$҄���,6'Y�'��.�*'���%����T;	���A��J�~	�ǮI|��N��9;�	�+9�tr���n�{Y�jʙ�d-�5B}��A�y=�8m����N��\��R�ŀ�2�R���+���G��p�8��7eFh&a�J�8��D�^�-c#�%����.pv�7��Հܖ �ps2x,Pͯ�;J��B%7F�\~��H�e�6�,�hm�������	^?�3�cx}��Ƥ�bA�%% �h�D!uӣ1��0(�4?E]�x:6q�]S+u��8ӄi�ec|�"�ښk�x�����-��<�@S;h4l�U�-�4�9#�0|
���n������A�����-%�]����h����d�d7bc�q@ى�6�ea2���Vu|�跴�@P��~��A�+�F�����,��lH�{���v'm�@���˘|T8{(��F�v��pլo�m'Q���+�$��ͽΥ	���nI/X��ou���T�AsLV'��zU�B�-�w{�0���D:��w#��h�c>S��vNK�UD��� 4ꌔ�Z=�v�l���5�	Qܯ�Am=�2JCl�D����O��`�
}��@|x�R&�����;��!���F��&P�4��&{�F{��uG���ˑ:�J_sʢ{׺�^�J���M&'�c�'�!�E��w5���Dr˵u��W_]Q�j���{tW���*s��Q��@6���凧$�po"���ل�������E#g���zf���I������?����p����}�)%.��^o����-�"�%W� ��y��=?@~�� ؍��Q���4SBe�������Ș"�y��4�T�%�<;�V>��v^��"���$�G߀)E*��/v��~
�a�%uO��I��rM��^e�*4�Lu�ٞ�q�� ���*:}x�oi�
������ŦG�q��zU���:i���C �u���8(=L�7%��`).m��������=ښ�ס��������9Ux���~�"q$�Ɔ�t�C��9�m�p'���r앢�_�}���+�[D����Q�� ��4p���}e�X!s�����9��o���\��=c�ֿH�AQ_^&���]7^ǌk�hɃy�[���
a�	�ڐ�2J���ي�5��M�[�~���BҢ� ��������ᰳP�(�=�6�dΦ�x˹�rC�B�{/i���`�@���qr�<�%:sz��ս���X��z�R"��ˉJ�F��X��}OA�%{��g	��n�?���V�_�yhў�PoI	��o7)��!���.��(/�L�����ɕf8��	��eƼ���0�1�����Q���~X�͋X�}�kR`>JwX�ێ�'}�@���e���)��17��{-��p<��P�R�7"�)�52��pm���3N�Ll>�B��6L5ؒ����ۦ��k3׎[6�aX#+�����	f_�VOLV�@�P�:�`V�ձ�z�!�m�l$2��d�qG�0�mۘ�zL(�,�d��v�fGk���h����<YK~S�S�����SA��d�ӑȢ$Y�D8���UΡS����ƽ�5T�͐�VT��Io�r R�YT�5g�F�{q�Y�)��R+�S�v�yc�~���`�'6��!/+�x�1<m���}��K�`d�;j��j�˳���u�@N��~ ༌��["r݅���{��EO�Z��\��$��2$J�ɵ]�X�ק,��}E%dΟ�f�<&\9�����T�m띪�z���r�|墘QF���v5<�O�J�SB�K�����(B���)U��������a��>ykD�Q�����r�̸@9�Ǧ0�jNB��d�D�C�N�P2�3\iwy�G�>#D��冾�vn�9k�%�ӄ���`����R��F������N���E��M.�� rQ	�lDx�����T-��~�v���ۃa�n��a��Y���װM�Y�Lp.Iײ�+�B�wf9��C�H�`k��A��B�H���3ףQ��f�G�#C?vf�j����0��N�!߫���K3�uV��9�!4%A�ɖ��(X�8��L��?�f��1�5%�C�&��d0��I��B��J��`U��Uar0�S�a�X��Q6��0Y;>Z��E`�9D�C2��vD?T��`�'Ė|Y���H&�L��{��o}�P_x�m����0�֘Qa"��B�ϕ�a�d�!��]-�$B˾�Ӆ�<ܼ?z��?l4N��,���jH���)���c{����^>00pZI#�9��on�lr�ҡ���~�B�y�x���$�M�;�=�%<'�2�&�Eiz�~�R9�i��6��ř���$SӲc\��D���Lr���<�<��qd�z�ڳQ�r�Lf*gy��-ڍ��u����:�Ec��-
�a��P-��>5_L�㊴�@z��G�}"�Df���X�#H\#
/Ij3_N(�:����=����tn��n�)��n�����X��� "��0 �{�{��;ǐ�� j�<�Z����8����3�S泲�Xiφ��z%�͜nQƲw�"2�`J1V��S)W�a3��r���B�#X\jkSjy2v91�F�&��D�;v�~��&_N?_'ZQ�n�=i6Y$�q!2�|���Q[��eĵ����!�)�����Y���C.��<V��Ge}�If[ѰF��աa��2����@3��ϟ�*s��t�˷	����^"/>[o/�3�����p����B���y�������'�P_m�bW��H�[QH���|�3���!~�6�zQ��߇��$0X��_F�=�����;�ȼ��+�̧��s�ϳ��-kU]s2k��Շw�F]�fI+pէ��3�-��A7&8@�;\>��$@b�B/'�a�|z����>h'��=R^m�#"oLD���g#�i	؊m	E�H=%2����`с�1��ޥ�/F.�n���3C�ƴ���IRMV��ш{^c2��&��1u�����m��Ϛ��W��XE2�ws�b�F�S���i�Z[I���ʇ&�P�7<����I�::̪u^��p���F�+$SR��l{��_$�?!.�}���]�I��V�4w�i�;�^yn��~Ң������F����~ȗ̬������zSã"پ���V!z/ I�}�tk&��}�����$t��SnM?�ӑ!^j�&�;`����=𘮣ě9��O��!����Q�Z��B��"��,��� F1e�|]�Pӻ���:_�{L�n�� T��Tod����V�ʛC���(
�4�� v�Win���� �*��*�'E ��ŮC+k�䳾�V�>1��ʆ:ڸi\���F�~j�+I��� /!a68T0��g�sf@%�Jz/c���Bn���!8&k{��U��␵CIg���Jm��P�[��vl3ƀ`mZ�I���ܨ���!	��hϦ�p�	��ۈ��9�Jqqqe?Ť�ƥ�;cN����,u
�,��<��qA���P�lgm��2J�i:���US��s�Ću;Z��U"�������Gs9G�����]��km>Ҋv�~�Eo�LdeU��\��M?4�S|M?���E�)p&���>������y]]�\^�)a��sս;m�����bEef-��b����鄅Μ9�nn���M�:�u.pO�"M��xn��^4����<�������h�bcG�_��Q��&�S g3<c��=�*���.7(�)½s�3?���-~J�<� w[�fB�J�),>���i���#��Y�[$�_<'���`*���('l��ZTѮ&��v��1O� /�lg����=�x�:��Q��A���gܧ�m٫�%D':B,�o�z퓋x�P�����kM^f�t3���"�g��l����F#KV����V��S<t��c�0cs�2��Ύ�i��d�Ͽ�.d=ڭ����<2�3�{Ƥ'�f!�p��R^h����BK���al�ۙ���f~Ì�͊f��Kˢ�yXe'�k�n͓C1��dzN�h���j��y�T�8k��C�M^N�{���F�Y�����(���j���\�nʽ\��^��QAf�)�у+5��W�����S��9*�� ������D�K\�R���qwHc�Њz���
 �$d3Y`	U��03�g��K�!(�Z�Q��ҲRO0���h�"N` ��f%!պ�PC���W���5"}O��q��`�NX`9z%�ggH�}��ٕV�b]���ox���.Qۇ���C%��s�F�	�ͮ��}�7�ͣ6�H�u b��A��G�U+K|0�J�65�E�y
���M:�{fMq[���	ͳ�gX#�c�Z��BNp�)D��b�vΝl�K�9.CX���~�E4������Mr�-�\�Q-��o��;a����o����yo�����S��
j�~�l��aU��na�}�	s�wPj@2u�1i��x1�<��z'�SV@ 0��x�+�;8Sx߃e�V-�h�����,=� =kIп[Un�6}�J0wD���t^��t�!���
C#1���n�=�*�{^͠	ExU�^9T�sЌ� �mWG��f��*�X���k|�A�P*��UL��E�.�1RU%���_��\��7�c31E˳��:����Gx��[�>�"i�s �~)���h����i�����m$ݾ:��)Z-Կ��.�Y�� m�%8���moWB"C�����aE��|N��$ ���'��s��u�H�E���<˽���׻*��|_�i�	�1D�vb�A�˼Q��c���g�e�>b�9$ Pe����e&��p���.��Nlޔ?i3���Ry�����	s/�D��h�QD�q��P�w�̸�X�Px�ZR����z�r�r�����ס�y���^VB��D��&�isR ĜQ_�N��oL~Q�K��d�}A�/��"���0D=.��3���s����9.3��V a<iI{䪯�UhV�Id�BGb��|��v��x�����hi��4l5Ql0Pfm�	�t#0�7/Us*��hU6�g0S��@�h��V��M�%��龎��ԩB�N��a��`�Yl�8���n2�"K.d�|�,��2���f�02����C.�]�-�R4��bjh���<��$�Y�i[_H2.W|	��E��/I�Q���ܲ?��Xw�4Qi)��!/e���(����%b=8�*�zK�B��4kݎ��=" �o��S˔Ҡ��r�X!ܳ=�i]/:@	x�v�(]J�X��c/MN�������;U ��o�ʫ���A-(��a���l���+˺k&��>�0l~N i(��P� �=�|�3���WAsW�OWtH�H[��]�%�2ѷ�e=�TQ���r�9͈.���WGPwu ��.!��fi�jw�<R`,�O��l\��[H+"&��bÙc%�qLm�&~I3{t�n��r��|�eb���T~B�L�k�g��+�y�ޞe���z|�[)� ��|c:��h�1���b��c㴥c 2��}�ɸS|V����P��-w�u`M�ԫ_B�ɸ�#y �0�(������{z�6�v�(qSp�x��ˎw���,�#��A�d!S��4�o��g(��֚
!��̐�<ؒ�t�K����RG&J�9�=ۨ�V��7u@@�z��~㋮#r@�?� ��{^���d��<��z�R&B��{c��p�G��������q�E�U�H��LKv��q�����M��W��hv���돬i-�oh���w�н��A�{�t�f�W�x��a�P>a���5g#6���P4K��/�h��C��YA�ۂ�S��K���0��?`��|ݒ)_�/�k�T�T�dϗ�8������q�ޝ3�P�R٫w�5���h��>��=�������J����J�P쁎���1��)���.�6�<$F!l0��|b���d�bP(nf�����CLL���VIV��uWzڷ旌�5��ܳ��<��C�vk8�Oɚ�V�a;�K��xN�,��T�Z|7����,ƫH�˥�S(������N?`jW�f!Az���1*u��2ڴfc>�/�a���\C�G��+�S���,]���Z������Ii<W�)xL��(�Rw��Fȼhဋ�<�<v�s��k���4�������
f*Cr�=�}��L�d1J�ܑjW���w�>F��n%a�@� ^��\��2��JF?葈��W�m.l�]!�q>�$y�j����=O��2!W�8���űQ=�2dQN��v����ä�p~>s�^�B�<+�	��l��^������6�(tNCjD�L�����9��֯Ob?%��D�X;��$����v�m�3�b�Q�+��@y[nw	��F=�%�t�L�#�B�Z�Z�X�5�T�b]�r}>É���+dsu����Z��0�
���k��\9�L9� 1��A.���0M�}F�(���Lv̥H@p�vyM�bi�i@vF@'������-��c-H=\��v��]qb^��� ]E��� � �W-P�P+���j@�A}4_ʎ�n�dW�&�r�(:�IA� rHh�'�� �?�Y
�zT�t5�D�m M�Ij�CY�a��-���&0�FnST�x�e�-m�a����ա$�t��\�z]�I�/��b�h����N�Mih�*�>:3=ԑOP�CT���:�w�rJ�����7"{ʭ=s/\?�$����rfp��m�����3,X�y��ʜs�3�}ԲL4Q��� w7���-�9>���u�ox8/��Ә��F��e�	���Y�I�
����]I���*�a��^��J�����(?j��<�*��G5��ؤC�^Q�_�;j�^����v�Q:)�-��T?#��!����b4��"ų+�]�N�E�1&u7��G>�H{)�C�sL:�y�\HO��u��1<zq����
k��`�_}%N-��*uc���`Vvi���j��<��ڑؕuJS�w�G�Ϗ�YM�KH��e��H������vR��X�4a}~����"J�B�<����la:�F].)��իcç�`�_��I}����9��_jeT��]%�pNFs�� r"i��TaR�M�EI��d��1�/�m�7�@LĆ�H�y�v��Od�,��?).�J+�1���%}�7/^�Pu��X�|�����V����Hɩ���1zz�q=F��� ���)�;'�o=w�8��H��wx�/��M���K��1�Ӆ��ӑߢw�#
�-7�?�;��EJg��"BI����yp>�U�.��B"���U����Y�Mj���N?I�8�qy�����9I�]mq�P�z��/�k�!�]w�m��;ǮFoU�xK!s��xH�V���~y��;u��m�&��̐<.c`pj'$��|�O�`K����NR\,�����sjѵ;�7J5���q>��V���"ޛ�]m�������c����z9��;�������鰣�݂Hf�Wr�s�Y1ްV>��|'�5�W�i;�n%r�&5�r�P�r_�[O�c��Z���bDr�IyZ��uƒ��d����)~!��=��N�'\W6�ƴ�ӂA�Wk���׉.��SD�8�O�}~v)�X���]�ՎJz�\
L-b�.,�c�r;�_E�/�o��`3�X�u��ވ�8����>�%6\G��Y�X�'~���=�+����+b#��o�C�������>�XL���� ��XB6����_!�-}[�?	�����y;�c|�`r<�)8@&�{��@)��%��WCz��:C9Ι��	�#�SC���'���|�R��Qp@��G��t�ϣ`}��>`k%࠵�\�?�6)+\��M�J�0��?Q�Q�'_��?oė*�O6��O�~��יae�Љ��Qp�֍�skZ1��ղ�o���5:�W�
�c��k��M4i��.`wz�I:xV�����t�y�d�ԷTUs&���/�Ǿ�*����y��W�1�H�N�%jp��S�<�/r;g�AN�2阖Im%Ԙ�U�|��ޏg�n5�o\�Əw��ϭ���|x!*��z�������H{R}Q��o�Nh�:�zU+-���n�#��?7H&oX���Ԛ�It��O�10� YA~��o�`�OCWu���^U�y��x�}�L��5�S�G�;��X,�-z5�w1T֑����cYm�w�7�!��d�['=�6n�Htm,�q����0H1�q���wT?A=CYTaǜ�(6�Tռ4��2+w���Z�<"���Se s�]�-H�&g����F%,���W�@��)�.) �# ^b*��|�%�⭶tY� u�
ȋı�pD���t�F���s�9�)��S�yw�P��w�4!v{T�H�ᐯA^Ж??���1�6H�;}���*sĨ�U��/�t�ǈ���Q=hR��D	��ՏR�%�o�Z;G�$�i����b2=�}U�%DH@`��� �����H?SkM�Cm�TP�F���V�R����m7�K������Nr�����qQ#_<��s˪�ʐN��,s�l�z�?j$ڻ%r�>���9G�ۈB��q���"�Wn�D�U�v:AtO J#f�&�G�Y��J����!���v����b�u�U4F�������:���ܣ�3��>m_��>B�k߹��p{jw$� ����ih�bW�����ծQ�ϝd\o��:�r�
�1���Jo������В,C���S`�P/��	d����V$��k��C��eW�n���ʩv�	����	��i@	7��p<�����/���l�A�a	)^���Oe�y_#Ͷ�7t�M�^Ԇ|�=�A�Cs*S�1"�$��L%�l��꜍��9CT���,"�I��1����S��$Ho�{¯-�ݑ�ȼ,�P�*D�P��+��A�:(,+r-�Z�W�h~Z��| �+��Rr�'��_%�V�-BļǴ-�8�8.bН @�,l@�+'���k�ʙ鷂=��y�n���1�y���v�F�{��M*���R��P��xO�3�&��/��:��´�9RҨ�#�lx���1{�dǰ�����;��,0�W!c�o0�n܏�
��D�n9����G��hft��B�'0�cɚ�#�"�y�Ȓ���/�MN�B��Р6��2��I=@~&��*���x 6~`y'��Dس�����$[-ƒ|��7 V�e[^ϗUg���-G
Ԇ�5}��s�v�1ec:q�'%d��-�4��`kq�V=��R*o\�ႁj��ڤLc�9��%���)�(s�[� ΅
z܎>�����+�.>�?v9��.Xqjcâ����u���� �(8��_��#:x�V�,d.�屡6���� Q�)O��7d6촡�r���C���#og�����${����s�)a����E���n.2=j>�P��q��rG&+����˘,���2����a�c�+==�U�2��\I��^y#�0\b9��F����sBj�@�� �W3���k��������";��K�hA�����hc��?zyC��J��:�*Xg�����X��0\���5����d��\��vK�9�7��7f�e?H�	(��Gj%���_�G�$��]�v!@qBi�g���s��-����i޾kU���y�!A�~~ާ��shJ����P�8&��:����dD_�[Kz���C�3�g`IT��hB
�v8?6۽q�ٞLg(IP���My)KY^:���~�w]diL���}�92X�*�[)����Q(6��� �|�s�C�h���1�>T����%FA}��0�l@�O��w��D�6�������\J�v�^[��G�<Ӹ�z���-3�(��s�G$��y���a#Jר�bƘ�0�!���Fs˹�!�f�Z��~���!�U|)xZ����~���PD��m�gv�c%��,+���3ԍ`A�\�_�C�(h�?���	��A����;�q,}SNE��К��3�7{�9o0�%x-�t�q���7D7�����ҥF,���b�;���!hJ�9�g�\�eWW`H�D�1ң�$�G}� �t�N�XR%�z}\�_Aˏ�A�Sט�Ze:�C�od��͇ �JB��\�"�=gx�J��B�uG�:@�sª���a��T�y%�P�Z�%!��P�;c��� ��s���[��:���4��x��͏��Dr����������-c4o�h���9{*��}[��::�v��L=8ޢ�E�Q)L�bż��i�-��*����.r}T�A,�b��"�e��u�U�D��A!c�n2�� ��e6S���/e��0>�UC��Ġ�x��L!����evu���� fD�3�+FJ*/��v��=S�s�o�����r/hu���y�8�"-�:��e˙��-@	�`�QO��$%n��s��aٹ��}z��b> ����3�?��%qy#C��6�O��� ��/�a�Y�Ź'N����ީȥml/��[�������^����g�82~��w��p�Lkt�/�?��Li2n�1�w�5&�������ق�fk���k�ҫWm�H=-����0A�A,[ۮ`�9���Vm�џ��#�m�||�c'1z����+�5u	��bRh#^?���j�\Ț��׼5�E7���{�IϜn,y=��k�~��b)��}��cE����(�!@T�����6�M(�C[2R��f�����~�w2(}!?vV�T��s���cŝ�p�"D��S����e]<�t��ƭ�r�8e�4�/]j�*K�a��jKaҾN���艈���|"�E0s��?�w�4Gkv��+5C���Nz��ar�k�J�=o�A���Mmg��ޗj�p	р0�nY�ⲝ+���O�{�N���qk���ac��eC�鞛�����S���V%��v���7�� ��U��\�|
Q0��o��;�'f2t,Y[u�e8p�ūU����>�/Z$z��X+d&�ض=|qp���p�e�_�.{����i[���)��b*���Q��9 VS�c_��B +�4���{�U�s�ֻ�O1�(�,�V[�kT��b���zP���r���i��"�]�*>�W)�KU�-X|�ӳ�a���X_f������&r���ի,�F��7ج0�4�D�Pӫ�@�$	�X��Ƅ�"Yl�'��	�|f��z�3��IJ�Af�ʣ�.2��H ΀yȱ:�1?��I!����)��|d6�ƫc�J���Z\�?kɼ����������3^�vzP�%�T�G�}���#T˼'�����~���M�-)q�������gX�������Y�W]*��~�K�ѳk*��w8J0�]�������&�Ln��y���[Z-��UI�`B��I�t�)��U��G�[�U׵
�q��H\�hU��2��ۆ�If,�����MI�Mw1��v�D>,�aB�\����Db� wh}��K�%|���E��>h���wDu����C$+�qB����C��F�"u�<�6?0����ј`�t�x����h��9��l�[p)JQ3�Yd�����5v��|a^�P�.g@�0��Z��`��k[�k���<E�ܯh��=]^��'���}���.U1T2G��p�`�8n%j���}ǩ�f�yP�~a|{�~	��	d�h�囲��2�ϛ_�ދփXW(��J;ҙĘi�3��]ϴ��k��eρ^̿�Y�>��� t�����V���ǌxA��63���X��g̓�[��<�"�V)e�2�� +K,���cJ0������>1c�]Q<jŘ-��Yg�C^���1�Euyp٭�ԧ���a�1Ĩ�WL�&�ms�@����q�`�S[�����?�
�C^0 q<��l���J��f�p(z����X<�n͢�tx���P�l�Zk]�&2
U�q���Y;Jc�l8
t�d�H>�Dw�0�~�3!��S?U	�\��B�
p�'_sLK�#M�e���Բ��d�?>V�z!K\h�}F�'��'bF�fVB<�++N�T��7�b�΁�@o�ˢ흳vSQ����$w�v]j�E��G�*�ݙ�k��[�t(�w�D����������2���T�T�����U��[�o�?��a�d4����@��J��+oF�m�i%W�3e�)Y�"��v7��׋�Y�f�@�t��I1Ro��7�J���$
eR��{�=�?��h(䙮�Y@�Oyye(0�Op�Nǎ!^����>�I�/C��w���z�����t�v�=\���`�1_˱�8�9��,kY��^B|+	��X�8mMxz7���1~� M��61`����:p���-D������
�o��BƂ����f.h�~�$�)g{`���H?6���V%;>��x�cl��	ڽE1'g �)�Kc��z�*7,9�|E5q6�u.������ַﰡ��I0�$��Eݱ��vL�Y��ٰ$Z&Bmדn�A�Y�-~���w Jn+��E��Qc��D�(�%�FuZ�I�C�#x9�U����$=�L�H���{�����5a}G�
-����g�d���>L?A��vf����ϣ���<�I���� Ezu _
� �>��>����7�Ȳ����3^Za%�Md~�2CZ���ug��Y�K��|�C����~��v�Z�)�i��j&e�>=:���� �ؿa������3c�\���}�n��G}Ob�.����e���V��I
��+,��o��T���7g�`�N��J�j^7�hxpg`��,�U�m��;�B>���*�v(#{�x�&���!��y�PR���n������j�_*�Z�g��/�Y~7X�E�n�7&���T��l۠l�l}��}�
a�қ-6�y����'V:�өD/��:	�h�?�[�g�ţ�W���P�^�ԟ���:?�n�^j������j�υ5���u<� �2)uY�,�Dࢀ���_e6*��" B��oNˮ�ʛ�]VnF4g�ⳛ�!Pg/x��$�x׻�Bn�ykȧy	�����k�7�UFrᦃpƾ��[��*��x5�2�I.�D�$�(���;���EjU�Ω�(��!	�bHr��M�]���V�C���H9� �T��AN���ܣ�+iw����r��Ӊ�=gykN�Z}��	@:Q���6�vL='#�<�����8Zص.e|;�Q�l�DJ�c��L����	vQ}.-y@d/إ��h��)YZ��J�sD#?JF��_i;��1���R�E���&g��"� K�5�����b�sߨ�I}�0q��y�$���\ٝ�x����"�*�9̰��i�a��f�$%�|BjW�������M�Fț{2�I�q}cC��D7so)°�b�^�vWȻL׽�F��.�&�s�_F�����a�	7ԁ���{(&�O�i;��T�w"�Oz>�yJ�p0Q',���N���ٯ��L���q�(��ڭzF��u�ch�V�7�*�C8���0�q�1y=*!s,�y4�6״:|�`q[�/c��AgK��Bல�6z�J�ӡ���ޠYG��1u�^\�$"}!���������Ի��;w`+�>}WG��э�Mr��_Ua���tU�8j���nl�v���FJ���M����^����td&���F��-����'��j�5�G�~qזN�p�vı�`�n)���� �.�A//M��gmD"����x�g-c������`ZT!q0��r�hX��p��YǮ _��ᮢ��	�
H.[{2%��R�ҡY�^8�q3��e���h*P?K6:��E�__)�ʗ���#>~I���g��?���i~f�ȶ��Ҕ�I����"��7`�,�)�`O�T�����^��ȕ6ʔ��7�Cq�o���:i�J��&���g�%��Ȍ�F/U��5gD�ɡ�m�