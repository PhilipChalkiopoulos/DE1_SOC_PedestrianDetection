��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z��4֬��9�A��;Un��Gh[�����<�#�L�-8�o����X0v�c�4��S�`U��� ik�{=�g]�C�+a
>kN}%]q�]���g��k���Y1��Ǟ�H� �a�C��O�m��ݒ�$��6�W~Zn��r�g�hc�n���,�+2��6�����Q�����ʘ��,&�����Q!�� >��*�Q�_tm��j�TVߎ��c? �E�^�X�������M�
6wbZP�i��|�ݑ����)K��*J|/:D����k5��p�|'����2#�[C|�����]�|i7Gj�́͑E���9�B�O!���P�t6�����A3o��Z<jML���.�6�?� �[I@xr�EJY���_Wx�{GN뤎�C�d�@8��,�X���"�F@���N%j�sJ7Z���4�����1��tP^�8�<�nS�µ��5Y��|#7*�Ä7��)c�H�+s~Oa~y2�V1t�H��~ D� a�?�>]�ā��줿o4,J�!	H(�s�����tT>� q�*���xo� Ց���z"*ѓ2�G��qn��uw� ޮÖ����m2#$)���P!:-G�?���G�e�Z�������WL$��%�>�x��
DCS[�GJ�J�(����4�K����n�SвK ��#������?l�7��/�C�g;�"��(̰�$~:���\iP�2�^���E{��w�~����������5a���� ����}��r��~� �"![��\ձ�Z�$'��z��f�Tz����'��x�m�B�*?�tu��ֻc���3F}��,]z����[�n���o�I ��>i٣��z�����u��f(��fO�+�N�,���D�=�J��WS���:��|~����J����.稝�k\���})a��z2ٻZ���"`s��8��V��m�.���gv]ђ/eI�= �&���Ήf<�?$�s��{�j��!�髁����E><��`Y�vl��^�ʧ��'za�=�m�K�0������i�f��,eB[JV�N�p�ڕt�B�ZXA���(���� �I�]U��@B�^�k$���G� �0�!&ư��ET��	͢�2g4(�ߐ |{����4�L��ɨ6މ��CǬP�	��!h0����E'�iM��騋y�1�UjU<�w�븬,��QN����Tekad���<7宰��xo�9��:] l�"�E�9�?��;MiW�Ӆ
1u�M*��x�X����Yx�;v�W��i�'^n>�J��ok~�2�!�b��Hγ	�`V���Z>�e?�;������m��׳Gw�/�r%�P��-!�IǢ e�h�U�:ǐN 4���D�\�#O�A�j���9�L�Л#t{>ET0���k����g���욺��P����j��p2a%;h��q��ו���yc����1��Q�A�;H�0�	��7�' �c�)mM������!�����`Q�*�م��y��`�]it�̡�QLHzT��{��ˍ ~�k+gw�٘�����R7r����;zϋ��mz�ѭ�;�%�g��J�V7\jl�]a���4������8��]� X�G��w���K���1#u-6{����e F_'9�(}	kk���a.썗��m�:z�H#0-b?7������A�+7�hR�J�#�h�=��ݮdc�1�R�}��´��rq��/�>��P��l"��,a�;�qK���o3�X	��u���d����P��eg�&/p�YSJaA��_�Y&�]H7j�G�J�f��Kj]��p�¤���>�ԧ�QJ�ORBhc����`)�<�j��ƚ/Eo�7��:_p7�S�{��&�������I���_�l�B�f�j�2�\�{@`�G"�{�ٹD�1|{]jas^�p�D;�JO�D�=�
�aV����[�A�l0�U���<�����`�A��^�M��r2	�9m,͈��My�m�GOZ�� Y�m%�#H�������t�A�M 0�W�6�[�jk}�@�T�{�[o�]"�#����AF��*Վ2�`���h3y�}`��(�C]�
��R?U�9�W&��[��q̶�����E����  �*��Ȱ^��p��Hf�����͏�����@��n�p�'Z�^%=
ͥ:���u!;D��u%�<@��5��RXpx'Q�M�E�w,S���V$A����`gdF�Rs!D��иY�F��h{��ڃ����N�)��n^û�����ud��U$B��s�&(��q��H:��y�{��_t;{C� l��(g	��:��{�E5&.�7L�Q�����pd���d"���4v�����.nt�{�19�v��
��i�b��<V�e��Z�+Ƀ8x��W��>Z����T�>"�����*c����Z�^��{�Km��s��_E����p>/k�K����"o���Ӥ:���`h��X�}Oh�K���7�_����"l���:˽����R,T>7��C	EF]+a�f�K�u���JK��H�Z��mM���C�P+�ї�5 R���Q��4Z��b�(8ebn���0�v��)�(�I^�z�j�a�*�b�zU�nݚ����u0/� ��oŵ:�JH��;t��"hz���EU�$ �]h��2���!��� ``9m��3i�gdy%sk�>�#SP ����KD���x�i�~B�y����Y6}یA�r߻��䒡rF�#x�l�>S׳�Qݗ<F靴T�u�87j@������m�K�t�g��=Y�n���-M&u����sY�dH�����/z���dKT_Kp	��Z)I����d���hU����Y�˗f/g�$�N=�A��Yu7�����S�:`xDdZ�X�Դ�$��@��A�y�L0�6NV���[2E�%&���9<��%FQ<��7�ũ��V�	f��(��]�q:N.:��2����<�d$�ӡ�c8P�W��h7�z���+��_([zK�y]�ӌ6�~m����G�˹�c�U!�+��3���:�=i �:�;)��~l�>՘P�j���h�V�ά��T[,��y��b��ƀY�j���?��2����L�㖍XP��a�ѓ�K��L�Fb���7Ϊယ�c1�Θw�����N^yб(�V�K�g����a����$΋7�T������J�p�6s�s�b�;�'�+��'�����h��?�n��Z�����}:��/3��a��J�4�4jc}�4����;{���r�O[{Eˀk��� ��E�P,�K��3���'��oT����̉�O8h�]� � S����Z	��-�&��GI��?���h�G��+1+t��_��z�cX��}`^Ǆg�lS�W!R�/������	_���Z����8��o�Ї@�(��#���P+L]:Ђ�p ��Xp}�>&SL9s� ��o��s�y���~�n#-��jA���S����X��}�u׫��ճ�����u�����F��_Q�ni����"���Sr�}u�����h��4�r��sCr�:_W�a�^�y�nK	�[q!
V���T����*�|�t��Bq��xY���p/Ly����!@��bC�;��#�>����|�BL� �9�N�R�Q�!�;����.��kqi+z�?���E�5��JLR�Ƚ�K&���{��'��	�^��|�ʲ9����A�����v��A�;T~;���(��Pt-��3!��;"�ʛ�� �89uj�_�ݫ�/����?[Ye�
���^v$La�$|�_3@=ڿ�(��3Z�I�/��
��M�5g}=W����>35�lI �)�[�l�S�,b��|���?�?ך������3�d2&y��}�v,�t�N>���=��e�`�'�uF��42�x��#�����Y���~�w�mu���F �Y��#JI2��6�-���[^�~�la���`�����U2�| ����H�\?�r��~�a���z<��CSgH��/��x����=°�u!�g�1͙LrE��������T�5j����"K�+�2�����pH'~x��Ι��n��,�LVJkWǁ��@��-��l��G7��ȗ�ce�6�/��+��ڦq��kqX��϶�6�<��+j�ij�&q���F�xt��T�=YIBKYd�6�J����+͓cP�qUY
o��1�'�g}}V~բ��]6�.]r�|p$�wW7��^����hvB7���ꃵʀ!�Zk���e/�����b)�j��L�gȐ��{^j���u�w���oO��Y�v�T�}����e�Bv�*��"�Pq�����8Uߖ�:'������d�_��{z��� P蟍KuUnPB��)��b��¸�]�ם%����X׍�]MO�FCk�0��FRˉ�e��-wc�U�Pv���3ź'��M�;c���1�-Fo��8^�/�P��ρ��4��umgs!P���مb����v�b�9r/.R�yҙP���_B�� [�o��k֜&9����ޜ��AT
����.	�NY�ǼIj���B	VO�,d99���Eb7<&=���AOM^����"���F���w���o^R1Z�^qvu �pR{s�o���!�.��#��<�bvY$�T���qPƅ*��]��cί����3�eI`K��_���Q�h�4E�9uO6�����॔z/��6��H�^�(o�NG�!"� <��p���%0��i��k ՜��7�˩ր׻ei�m4%�@V�M���S������WS=�1�ToVRuȝ7U�*2�����2y(�&����+;��8�!�(�v��Ȥ�$�-m���}I��V��\�D�&��V�6/�:%��d�Cɜ?�v&��#G9�bw�f" 3l�5a�6)<-ܟ��+��B(s6Q�fU���|�3�;v2!���M���6[�"떶T��<�}@&0��X3�.���6�-�t��A��I�b���p9ܵk�mv8�V���|��^yY-��5隷%t���*B�TY,���>�` ��O�2�usE@N��5��nϋ����Q"�������Ho�;�uK�MW��T���)w[�]��b�N�=#��8wc�ӿ����gHQ�F��*Xє,��v�f8c]@oie؅�ގI$Rj��D� �*�^�O��<���[�K�W/%�I�O-���,Ż��a�p9���MJ�M閳?���G��S=Y�v��$Q�>Ftm0ϑ)l}�m����J�3bw	�s��bE��O\rL�&�,[��v�o�����ʎ�U ��J�5�uL���y�P�f>��q��Gl���iݿ5*..�^3����[���Z�j S�D�R�,����\;f�
$�*)q���'x�
�RL������W�n ��O���zmE�s���ɗEI�\Ϝt���Y[R��ʓ���)P�F�ܧ+�h�#HAf�ld�fU����i&H�OTY��{���V�G�~LR�$�`�<Ab�q��:�G�Z��艆��NΗҁ�,����G!��u�kQ+��B/B��'�%Ѫo���	X��uu�.���.h:?(�C:�ӎ��WaJ��o��R�px����v�ݺ��u��HJpQ��������Pa��u����,�{�����rJ����O���ȫ+0~�\��M���'EH)E�2���W 5�|��^��94|b\�/�pe����}�z������.Uc�=��I��W��U�M*��.���a��p�ͳG.:���"��t��{��C+&r҂�;��g���VϹ��8�$ND?�I`˂�0��
A"�%Ц��E��!3Ơ9�^`��u�$��f,R�"�|+����YU����,��S�6�034"#�nAj��[��#�)�����i�i4ϭ_���V�o_�]Wϔ��ƒQ~ �Yn�LQJ{���i���-�P�֪ԪW�Q����b��Չ����)A���ZR��:rik�/�C��&����3��r],�n}z{���6��|SN��*����G"�W�R���s���w��Hܒ&#P�k"ύOfgqˏ)`��z,Om����y��ސ���7	��O�@�Dn�5ˎ�U��x�����渠#�Qq&�K(
NR�{�<K��6NT�_����+��uu0�P�;��̏��mʥ�@���SN�%��(�DԠf��Z�K�2��f���d��a����s�7==N F�Y7^�t5u6bjqC�K�D�c��A1��+9��m�C���r藧)F
0kr�|(|]���ޟn��������;�}�&s�=0�,�qi��u=(��"<؊�@r	�-�IRn}K�㲘����!�Sa���_I���)q���q��}
���e���Y��J^���+�k_�q)Sv�
�J�tr!ȉU�.m@���}�7a~(oA�h���:d�J3!FQ�wǍ6��b��Yq��5��.���W�z
׸�CF	���Λ�"S��`�S1�U�������� )�f�;�u!�E^�辖8���\�e�6�u&��ҧ��x��S�����}*��(�GVkmo��P���U�����I9�oW
V�LfZ��=��� �)�&�r����p���K��y�va�5=��T7�)���h�
���l�c	Ҳ�/q���(��c�2��,x4fd�
�P�}��Ȓ�ƹ]�F�<�����K��X�~R�i��� 512n� ��D�~n2x�W����Ov�Ԇr���˖�h�#�<�"o$��!�h��:��UU��~v%�0^[���;�<���"���!y]sh�t0"����I�n*�$	"�H���?�H�"��P�&Y�K��Y�-�,Ĵ���+Ę��U�Q�5ja�V`�h@�h�89>9(h�D�B�:@�G9~v���z�}�~V�6��f�7�1��-C�g����(��>��A�$���7F�h�+i&�a�?b�=ۖ9���8`/\�69I;�1��P�Ջ�+���o^#���g��ޫ2�)�av��:����+3�Y�{��4�n� ���^pi���4�B�k�9�<}���ҽ�n-C}F�%n�S�$�n�������@c�H�4�
;dbrw����%2^$.���u7��F̄s�����Sty�z2��џ=�<���Dx��h��ӽ6���� ^�Zl� h��t�Q�|�?kD�����g��2�]�����/����y��ɋ����?��A�&��F�8�!6�<��W��,=��h�LX��%��б"Ӗ��6��f��~�O �ۍ`2'T���ۤ������ɉ
U�	���u�����H�L&��p债7�A�����kq�29.�	,�ʅ;��e��_��Ͱ"��2v�R�ctΚ�tY�8)Ɛ��E�~��KR��N6}o��)5c�G՝�v�)�� y&5�Z\z1�Kbq�AC�'�����B*����>��0�>w-OH��	��X�k���HϲR���*c�V`� �"eeV��,��0�yo��$qe��*�YU�$�?W������֝����qLe)L43�bh/�a2Y��T�@_z��� �Dѭ5d2sd�o����Ox��|�Q�d��UP�.Z�D�UδB�7\v�߭SapEL��-_��Jb��ʽy��,�-�.
zb/�+IW"�b����Zh鱙���-f@'������#%���+��������£f"��Z�l)W�{n|^�3�ɭ�O	�]�,�1�4���F�7�s�`_��-�}П�_/��B7	s��ݩ��H�eRB��H�{5�#B�0�ƻ�u��HO��2����$�Y1���*��
`��W��>g���R��<]s�[�&�V�R#�T@\r���j+��t��wo���c��n���o��8���TЬi)I<�%�[/���'(�ȿǎM����,����|���˸�X��l�|0;(�
B+p�Խ��q3o9���zi!��:��N�y�DǺ���� ��T�����m�;�p�Ef��Q6߽�T����0MT�P�ЧT���y4.��b2�4�r�����q7M ���A�b���Co,�PZ�&�qbb�>|4�>)e��&kY�I�tg��b�玳����W�׉��H7ztFFQVvj���B�;b�!��a�����1Oʯ�\��%�}$\GH3��Ved ld��l3����eD��ad(ȹC��O�z"��_`�qbi��v[�+�Hy,�S�Fy��?-N��a������*��a����\�!N���ЂC���4ZT4Np
���p2�	�3����>8o�b���\~�
v	R(#N��8�n��a�aq��7urkM��J��xf,�Xټ�Eh���N�w�n����K

��M!I���!o�e���2�e�/ TQ;�` '$Ԉ\pׯ��}������T�KzZo��Yl䭗�*��VFl�z�/�5��=Q�d
<�ޝlC��(L���7=�Fr᳴�wF/�p�)|��_O�H]���*�%rxs:�1����7��Pl�c7c_�#�wA�zY�.c�?)B-��[IV}���0VgM<��<Z"��Y��G��}�K~�֢�Z�����+.��O���S��h����NILj��m�`R\��3E�&+�����V���M�V�޴Z!�-%~�O;�g!�,�oM0	��(1eSpP�e���A���
u�6�?籏��Ƕܞ*�Z��E��LS
}G�$=���0�'+2�@���I6[��#�9M�wΫ&b�����Uy�ZW���⾭�6{�W}t�l#�,4
�s���f��.�[iȯ��9��jم&BP�Q*��X.>��Ʋ��9g:B���@���KB/�Q�c�o|�/��p�"0{�����v�M8�F&}v��^����0����t�38�NW�"k�!sX�R��pÓ0��+2�ճSU_(��������˯:O�Y�F�N��}��W��4��àǊ���� c��}��n���,R��u
�.�1�x���{�P�cQ_fʛ��������G�d��f��	ɹ���d	�����2]�!©�9�2�u�j��Ț��6�\�=z���91�-l�l� UZ��e��|��p'7�/���d���Ѣ���d�m�~X����IS'
��@Ҽ�� �O��}ղc�A�*i-9�Y��s g���1/�u�V�`>{`�ubX��]�F^����^v���sD(d	�V�^�mO���oۗ��Pz�ꆯ�fh����Ͱˎ���w��v�m߆&Fnj`��������[9�Aꨁ;��>xR�'"�+��@��C��e�9LGC������%Wܦ�==Z�q��ܿ�zb��Kt��G6�!�������U��m�N��箳88Dd�cf������UC�����v"3��Nn`d�5��t�»#[�Lٌ�����O���ŏ挿��S@bg��I)������ 8`�e5�\��8�Q�m|Y���s�TG�����^�e�F
������泔��'�E��T�lÃCy#�%_b7�$��<M_9 2y�����+'w��ͯ	_3=p���>r�+��eMO��D�.ʵ2����4/��.T�O��#6��X�R�A�?Q^QF�"b=�?3RWv��gױS�6c�h����:��g�r�y?�C���"�$r�[�&�_=�ΤƮ'������kw���P�$��,ƞ�	j
Z����Eg�����f����m�8e��p��)Fv�8�k��M{�����*0R�J)ol��@�G�#�1xY���/���+Kt|䆥��+�e�E�Q�h�?�T�.���)��,ҐHye+�%*�^(����ߩn���ȟ/2T�k�U�,���L�$�M�`��ν����@�ȅ��e��dٺ X�3����
żu�`惺��/�vmj� �g�,�#W���CV`Fl���}����6\�l�g�iB� ���2�%���-㾨�?;��P���]�]�~{��a>��'K[�wl�EK\W�雤��-T������؉4r��g���޶��������j<��j,��1�e��O'3Q-���诌"�]T>��0�����ja�?D�G�0y���KI�+�&?Q2I��, m����u��I_�/Ĝ(\�fa�<{F:����gQ�'�5G�9Z_=�~�C��5�����x�	o_�=�C/�`JL�&7�� >hR]�"*���42	 5/�;g�a�<����5�wQ�@e�#����w��%��4��Gs.�n�+�W���4����a�P��<ُ�V�&hQ~��� �s3Cw�i��T�����Ŕ}�����G�;C|�vq��{P���m��4
i\1�ۘ���j�AW�mz��\��$D��m�`8^.s�����"iJ�-�uK�W;%���e�R	b�q�AO����U�k��Qt>A�+�(�ȃ��e3%v���ȝ�I����ԩU��;���A��\6�r"l�x#���3A�7�4^�;�̚�j3y��A��T���B�Q%|��'�y�
�e!M�J;5���E&�k�g+�<!�����~E�Lk޾t,"Ͷ-"��L�%)n�>��U������J]S���5����*ӹ����ȧ�E��if�[����(�8Y-�_�7�,]�~&�v�P��/E���� ɭ#p��w�RZ�"�5<Uw�;�$�L�}��W��/:<%5tڽ ��sEn�՘��RH�㨎1��l�gQ�ET�Y&坼�Ŕ��u�>�yCw"���!�t�Z7�KyxR��4v�����x\w 4�Ǜ��k���ܪg�ER�Cs}��,��"��r �)y��Q6��E=QcŁ8�&���#��2wt�$
{���gnm����M	Lry���i��{��vFO���ҍ�%�~#��X)�o�4�o�����Ӗv0�	`�^OjfЪ�߬����턜/�F�Yy��f�C�1^+KH(b]]�DQp��EH�)�Ũ����Zyt���V�,����?k��@~[��H��%8TUB��Қ#(JR�T���j~GR�^���ޡ¶��j�&����,�c
�����Q������d�k0�4���b��iC?�/�b�%A⣔��Utk+GS�qb]�Ձ��Y�����)$T՞�/̢>����6t}X�τ�$������;إϱHoWALǻ4/zF��V��h3bl����Tu�G����̙���e!�N�K�Au��9,ޚj�?�4�
\2������ 	��
�6�>*5�~���&d=�ghv-���f�Y5�B����#g@Dy#��tH�a�d?��@zb!�L�:�Z=��%��z)�$_��pqV�a�;Xmv^�j�gR����tT�����w9̼a�F���d	��T))!`��!a$�W:��u!��,ɖ�A�ɸ�b��įY��b
ЊK��A?ъ�$8!~0�t��;��"��K]��"��l�s�nAB�Mܰ�N�)�h��r�����������,��'^K��F��]}bff)��AȀ�o��V��P?��zy��	r�Q��J��e�����L�pL�M��֎rP��#���h4�n���}�+)��6�ȼ�zU���3��dx�+��C�W����?�4~҆6X��/��b�j�i`����,~6EЌí��@y@���?���牦�U�o[���$���%�'�k��ӑ0���q��C��5��uٚi�f�I|�K �9َ���1�B*����dX�Q���b[��y	���]t��Lj�E����i����y��������<�dG��4�h&���)�0��=�����y���� ��Lu�چ8,#�1W������} �)�	őG���������"8��Ʈ���}��J��({���t�y� UtSɹv�Q��!�^�E��ۨ�5#F�;��\��ͳ܋0�G;6�����s����,f��z4�T���?&r*�pu�8*4��g�*�19�uc'��>E��u�j�2i]�����\�����if6ٻ,�Z��!�f�����g��Uh@o��V��UHs�V}�e]�7+=v��W�4��L��vK51��\ "}���b����!��Y�/v R�)H�S;�O)�o	T�Z/_Rɂ�3r��\�,W��݂r�p�hyضVP��� �?�6_�Aa:�\�X@{��x&!��U���B�p�=?B��`�b[֙�R���yû�az��`�d�'�n�ɵu�������/v �s̼�{��<l(��:�������k�l�<T{�D���ͧ�#��|�%�8>Y�h5��%��?��XL=M5�/R�5�Q1�oup݋w����C��P�G��Y��5ݪ��u����+�gQ�+���'KlA�iLjg׹�X�w�9e�\�ռ�n��A9m����K�n���z@��Sz����6Ө�x���U
9��vMr1Y�NF�%������<��D��7���s4��oI�M��zGC�<u���f��7�H�U{ oA��m���������V�yB��II�Sm�S��YC�i%���K<X��yҁG�t�;E��N�'xh Kv��z��p�퐰"_��'N�a*I�'�a�5PIKY#	%�(��άR&�~�쑶���I�d-�I������Bt4�J,��	UD-����\�E��ŘR���~�Z�#OqO��X��~97���q��*�$JJ�E�d{�0e�)y�i������74��u��A13&�&�@H*�L�2"6-hy��n����F�O�<l���z�Qr%��0����9���]<�܇�&�m�0��6�@�NM���#W.��[T�O����2�D��*���'�>�I��CJPr}M���j:g�wк�)P�%�y������� D�9u�ZG�(����� ���\�q!m>�3�0o�<�0�*A�ĉ���Ы��%��Z���Q�YH`3-r��N��W,���K�x�l��&r��yF��8��ײ��*��O�Ui� P�
6����"y ��Ԭ�<M�g�[�)�<k;9��"d����3�]���RX0�]�y��K��K��S��^�n>u��G4��9g#����h|�i��8�j�!�}_�!��.�����e^Y$���/�å�H���\~��6_=���zar�	ǈG�a�+t�uXEutJ�B#�)��)ZC ��+U�v�f��%�E�5rd�-m��O�4ö�\w���`�p@)��L�&
E�
�&Sƴ�æ�^��CB�;%z�<�y�/�����[�7��س�CQ������A�S���!�-HS��Y�9T� ���뎧� �Sx��Ű��
��v.�T�k�7�$�Ql�Yp;E�[��� �υ,	_���Z�y��4�c���igD�Dp�J��ۦ�M��	�	�=:�7Φ�o�g[�J.u��វߛ�ie��v�?p�����b��ٱq[EוA���>x�̚����݆A��&�w)�:OYP�^Q̫9ձR�-�rζb����(њ�u�� i瘟l�=�ҠC�1���>�j��b( �9����f�Ku�GzK�]�|�4�]+��-)��$8��q���j�/�0}��z�e�&:f/�C�0\l�|�,�JI��S,[�.N1꟏�F_��,����&��d6�,�R7��8��8ն����%�G�X���
ff�����R�'�5��~1i��$3���V�����l.
��p�ʘ���6X�z��g}���2O��~5	��a�����j�W���"�Y���������yfj�:oInc0�j~��j�AHꪶ'��|��q�_>����p� ���9IA�O�,9��fO	e� �{��a���� Ep�
�&�3&�T(�p��#��J����c�������0݄ދj�m�;ЮTAVj�Bqy��Z�}u>�G��Vz��ظ��l��(�>�驳rAx�̡0 z綸FVf��+$�c�+c�yoa`v��D5F��P@@O
2�/�sأ�9	�x�L�./��C�1g����,?�v@��z<�Q$ט��WRڔ�Ge���<M��]n����bs�Z�"?>�ڶeU?�2��$@�/�>f�^������[XLa������U	룖E�5
�2��&�Z�^�8��Zt��Y�je��ixr;�X��▪�W_lFWɍ����A�����>D��l�{b�vM򸜄O�̾'��&š̒�T@�M7���3dn��-�4<��y�4߿Y��Lj5�? z�n�Ȟ@�8B��,ٶ�]M~���RN��t� �02��Kk�j�/yd�Ohj>�8y$������ �6������ws���Az����5�Ź��i��ӚiQƫ�~��,���3�E�����t<xI{��Y�^B۾�ר6K���mӕ��N�^X�Em��D>zu7�}��ؼ�%�J	�H����3e����̧�{���KY�Y(l{iX �E���
�S�f\\��@��up��T!��X���)[�ngiQ5�<����6�C׋���jq$�(m%8|z�$'u2��Q��r�<�����a]����#�R_/��a�˃����R�&�eJzux���:�?����'��tc���j������5v�ĸT��
�v�A"D���V�X*ϣ�±@�U�O�%�y)@��g�?�����$����,�
1sk�b{s�5�j�M"%Z�1&l��J�N5ěr�d�W|�jE�j	̄?�R�I�#��J�!�G#���UTf{9�1L�C7�~p^��ۓNJ����v"r�(bK�@(
j�`o*r����K[�j����qb}k�w�����QR��"��$�8���$z�hL2()E� � �˲^���ˑ�D3nj�e��g�A @N}�'�IYy��C��G��t8`�Nz6����KKrj_��VZ�����g��l�Q=�y�%��@d�+�G���j�y����?	�[S�M��N�P����86Kq����m�X��C.[N�M++\�>n�m/���Ӷ-�ɡ�/�KHb��_�:E xZ"D@�9�,����*j�iqO ���������ޝV�$�u(嵮%s~�����S�u�S*І4� ��3��˗���1����D]�ǘ��(��o%����p���1�~���T�����-'k�;g@?5����2�x.�<�T���L������/�Ws�Q*�30���F2�+|��B��f	��A
`�!R���0Q���@�w�QE����}�FRGDY3�)b0�>9�ݾV��!�����EK�c�Q���d(p�^S߉,&�7ݭ�X� ��X�����*�NCɒ�a��X㝛<1�ƛi��<�bl
 Y\����rM�
��7ٔ9n$xc|7�/%,HZR��E���d�^�k���ԯP�
Ք���Yo�8��Q�E4T�2��@-��k��i����?��ǒS�	q���Q+�I	�)"#��m`� ͟z�S�x���`�}eW{
׀1F�I��S�5톕��f�Vp�'���S=�~*>�W�ْ�b��k�-L����N��S��7�9�M�T9�iKc���\�����F�/+�U����,��}�M-��"wCK�w6� c�e��W��� Q�w�n�A�����%��'�{Nk�G=>*��>�)vTW
�=���R����mi���Wd7�Bwmf��93��@�ɺ����vF7��ADCg��(���-�aI���ܸ�Z�:h�����H�q�( ��~ ��%Aj����U]wL%����f3��p�c�S=9�{|�ޤp#7>�u[˦�o����d$�Q�{k��I��t�au~��w��-���5��H��;��0�a��2���V��}�ù�o�@��r��B�छ�1�� �K�=`十�B�IO�n� ���i�\�5w�U��晩Iu�,1�Vp��*^`2�d�pX����60����/"l���*��?5��*M�A����G$C���Y&�U���OxM .}�?��K���s�g�$p��9��Lv
#�qq��{.�a�3q�#&��v�+�/\ұ]<���*��P�-o��ӍH-i�{��A��=����H�h�;~�D�Q�^��P<�����9Q7��镽Vܘ��7�����PK���bݕ�J1���(8��\gIZ��W,�ѢKMr�8*ɀʫoA�<�6h%�'���?���470�wk���+��?�EΫ>]@��gW+i�=�g�7���y�<�I��j:��m��@�a]j��g� P����UFF	��ݚ�?9���d��o�Z�\���om�P�5�<� 7�@zqhEO���g?�XT=�L�|Ù�R�����G�5?��۹#q����"���[����؇��nq�CHr��N8��hcW�?����)���q�K#~������S��ź�����^�y�L��O�\��}�F������}1�r��ǵ�L���.�X����ñ���p��F����@����� C$�n���2Kɳ��;�w�/2UM�!s���=~�2d3��lC����m�K�2���1{��/4߶[���M$S��#D�~9���8����7�A�VMh�+ g��s�O���
���^����p]�r�S��+��m��6����e"Q��p��W>�K�<���2�zu\��DD#�Ka�.��C�Q�P��K��׃��F_Y���I�k�9��-��j#%PR!f��������g~�!M���W�hC�,���e�/=C��[p��S�u��k
ȼql}���ŉ��Sе;d�6G~�lL\�9�i�c�y��k� �c�ɺ�:��t26���b���}�,e�|��+�۳���Z��,�%�wY/��Yg젝&(�>���V)��w쥭���4�b_|/f�5٧�>D���Nt}���6#��U�l&� �3�U}��d���EU���7�F%�d�jGh�+�}vc\����F:��Z��Dt���F��U�d��Ց]��t�	���Q���ă��G�?_`�D[7p�̗zO�U�<y.jyh��@k��j�
��טbʠ�3"Sk�k��b<�A^l(����a��*�K�{f:� >c)��V����a1Ǿ�T";q����"J��_��2���	����xr�j���ߓ�L'MI��w
}
��h�M$*Z�s�?��*0��&��y����� ^̆�����^^�r¨X��y(��,�cݧ*��tL;\l��=�C��o>	�EJ������������f9Kf�48��h�`�S#^+�=>���,��l�Krt��+-�e�;G���f���PU�б+�3��O��z&��}��<*$&���1������^��vf��$[6L|k��9J�$@�+n�<���ר��x7��Ĥ���%��؈$N0}�#�	e��Ϊ�R�͘AoN�>�cʱt���B�ɪ9�]��uԼ&��:�e��Qa'J-��v�zऺ\4{�bw�U?zAI�XK�b`ґj�~�9�7�����-���S�"�g�OP`�]�S����f}0�qM�0@CM�Р_I(~i&�QC�I��;`�[ɟ򙣺��q�t�9Q����H�Ǉ�K�h�B?A|�&�����$�a���
����"�\G�3�{%*J��鞏G�҅w
J�({���.f������6��d'9.�7s��/-zz�L���ީ,��pǰ���[�G�n,���*t���8��*���r��^Ý ,M���б\7x�HUtgI��.6��X�u#��ʐ�=�p㧟�
��+ I��g�������@�c&�j�����]�d����ip�U���-0qRF�cĦR]�0��qT|�9�F��O7��(n7�V��cW
k$2�L'7J�	�����"�B����]UL3��.#<��y�r��i��ɪ7W��ԺP�g# 2�u��PddUS�]մ�c7��rz�A���c�rH�R͘�l���ȴN���%�����b�Ej� e7o�%F��m+w<VA�>��7�h��*M6��,�ޫY���N>�j�&�k���A��ۥ�ޔ�����ғ��='+�3w����G2�nUC��C�s ��#3��(>��A�5U��~T����5Q�`	ծ]��dȹ.L�e>�(n���3׫0eDM���Y�{Ȟ���?+��[�Qw�Hs�J2�hB$�޸?~�^ѭ��mrtV����{����h1�ͣ�F����Y�=����Ve�XG �ߔ"R��(�HJ��lr�e�|��ev�74�\�X�����gȬ�F���~��I�RÓ��
h:�tBȹ�}�fh�e�~>Qt�����$�������2N���)�!K%dgB8� �u���N��z�Y����D�Ya\/J'E׿���h��
�Gֻ �[�x��!����3�*
a���E�Oh��E���j�>�{zx�i��2�dDQ�w|2֗K��k�.凋�<P�>u~�$sr�@��5i�S�`x��T81�~�ue����z�����^Pf�z���3#Op!�o�ᑲ��y��>< ��-���gQmDL�t�C��F��P�C2����������3���9��Q�|��7��ȏ�߅P���Gh���R07��q��wF�����:F�<��Ր]Vӕ0JJ�+���~K7���P�Ў���\�w~ `W�+)��\�#F��`�Y0�
0�YI�@
K'�	%�0�(�RP������3C�~IS�j�WlH`@���ɻʲ�o��qW|A�O�n���'}�8�"�@]<�神֎��
���#���Z�+&���?�_�~���#�u����2�L���m]�|B6I�;o>\�&��,�z���%ݛUJl�8���B;�)B��ja��UU�IM񮦀!��tc�q�M�.@�P,Q��p���7C������"���sI+c�:�a:k4����N��Ī<��E@�������� r��O�[��&@�a��Z^������U����2����zUA.�W�NB���e�׈భ�$�Q/���� ����Zc�s���B�ˡH,~WV��{�n�.y!�&t_\\��W$�����1�Y����@]�&G?�=Ӈ����3R�)8$������4N�&=�c�������q;vI��F�w�!u(#�0J�g�I��<u�����앸n�g��a;s'�Z��]��v3�z��W��m�Fy�O�xl��{�S���_�fub�&�g��Zz�y�oC[����hlS��������P�!�kMw�dT(>��g(dm�<|���e>��]�sw�
�0#Ư���f��J"<`@Z����,��v\$��;�+�e�~r�;r��G�1G�C߉�T��G�c�$����八_�h��_���W�F%�h#�p��u �j��%� ���ܙ�U��+7'��'���jI6H��\k��mZ��L��39��G�����Ww�� �D/W�~%��*},v�Z-wȯ�|\� ��%g��RT�����G��!���7��k`����� n�� |a�pf2����w��袄:���\�␻Isb�
���)�e|�!Ź��wtt0�4��iC!���=��A�7i��C��Ί<�xq�5Yw����1���\�U��-zӑ軂eD��3�焿#Y��!�%�k��+��=�rt���!�j��dmQUf�H�),�����ZZ�rI	�|5yn|�W<�Z��bY!��f��l��[n[�I���fh����a�^����0���J����7h�]A'KI-�5q�=:��o/k`���*�y��v�Zh�ДD.�`��s��B��2������I�7��#��(=҇�v�6�X����1+��>�`˸��|Yj�P��*�\��� �����Y1hp�]���櫵:2In�ј�|��ME��)�Y��Xw�QZa���		��j�x����W��$,oJ��Yb�SA?:��%(ϘÂ�̭��(q���l�����6ec�gX]6�����-Ev�ܒ�� R*�&`Zh�"ܺ���i�����[b5�TIeio1�Ҁ��]�a�������F�Hgn���:FɁ�ĥ��r]p�
��z�AK���C���b����q��.���dDL�cp���LFq�q���q.�ݽVNW��W���� 2��ίׅ�+¸c���״�nOR��s��[���M��phwq��n�)�!���8D��H�f�Khg�N�W�4��B��"�HUT�F0Z=����*C�NM�_�m+�4!��:l�ǩ̍�B�z���`��Et�D�TIUNDżɁj-Zw��䦻��,I�-L4O&_���Xe�v$J�?`�Y5��b���hR��&a��bM�3eʢ	{f4:@𷛨XȎ!J<ț�c�h`tdZ}�rʨ��%@�l	�p�1�~�����d����6�*%�>��$�fe�K�T~���Q+�yM�߃�t9D-Єqi��E	��շcR�&� g��%�&� #����+��9&�{$' ��{X���q���I�0�i�����	�b<��[���ʨ��A*!ק�w_&�mٽ��ek�f�;�qN�SQ3�ѫl��;d��x�ޕ]B_�ą�\'�+=��~��]8�;�?��9�U�';-�}4F�]�SKv�'5��T�_��������v��9�3��1=�7v.�C�y� ����v��kD�i�Q�ɡ'�慏��Ӆ�N$j�J�	�ű�K���9���!y��"
��,O��,=	���lN��E��%���Wǖ��H����v��H��r%ik��w�|���h�}����yX}-�l1^���Q��mCM2}Qw!�2l��|zjy��S�Ì~^dP��,�5�����۰�x��!?G���"�oݤC<�>�R��<�	�R�O.��@
+�=Z��|YÝ�RB���*`���Md<Z�Z0��@_#�2s/<Dq�* V�:	�<���e�1S�_XV}I�lʲA�ă����q5��Rd몪�G/����& "�EW{�0k�racGq���7�q���2Nyk�}�j�fk*��,c)��[L�����!�Qe���c�DW�%N=	ʥ�VUE ���\�����P���2Y�c,J��R����G"(�X��`�&�H��q��<7��ꅨ-�����1��Ry28�������|�hD^.���Q�P��/k�'��l�{�".	]�4k]T�ŶT���%-�6�K�9�{3�Ƨm�H��ҍNk�'#`��f���1�c��/)~��.==�a��ą��I�{n���mNy�fU�}���jةɱ��C��H���+�T ꞈ9��|ț��-��B�*:z�l��\p	L2�B]��ED
Hx� m�X1��6����r�Lċ_bsÃ[���3��l�U�"����g9n��Kۿ��m��U`~,+��>_�
0�ه��vh�>WCN�j�<Q���{�L��D��y��+���b�U�6�\��5��Q �����!�>�������|;E�)�Q����UmB#��X�<�>���S����]� ���+����Ij��	&��H*����9�<jI�B[U��)<f=h8M��-�]�e�����i����Q2	�lJ�ɖA�P_ƈ��?���ub,JH�U�Mw����H�J5�7�)�Ƀ�Z<��N�
׺�{��i��pĹ��۬
�H|�o�[Mno���-c��	a�;z݊�z�z�?���(�6�w�S/^�8��k���-h�H�/h��ǂ�t�Tah����sj�dM��S�,��+�0o�GK�N;qex�@%{�ﳨ��fI�",p�[ji���`S����t��:B j���/�}W�,�a2^}�I��Iq��'s�,񽻅1���p�)F���@~�>���ls�[B�g��f�S�,�mp� ��|�#�G�7���䢱��"�!Ceeh!��DMd�&�3�U��r/���S�(�}��v8�ឧ-�-��	d���K�Lfu�3U��.-c�b�K���j�6�>Y�yS.O���f���J(0%�w�<�"�\Eԗ�3�w�j����#��`=ٞZ�̿����R�t� �6����*P߫c�oU,�G�Mq�S!�]SV��[>�ֳ�0N'�=��qE#>\$��e_,zt ���5bx�qcuCX�#��0y����x�vo�!�ф�W�K���N:C���!t��E����c�o��%��r�����;3e��l�
�f����,"X���_�^>��g�4���-��>��o�����Í�Z�ڟ�O�7]��;]Y�MQ�P�$y���ب��+׶����cǔ)}�������G(䖓G�兔�<_���o���)�PL��'�h��%��� ��0X#����2U�ScZt��L����R���,���N�IH��%&;8���6Ԙt�-�,��R�wm��o�S���2�6�7��c9[?��rx�-+E�$�3O�;{�!�;̏4�&�%S�I��>�&$	Q8��k~�ٱ�|��ʈ�m�Seo�6�W�����wް�ؙ�6C�%�=�7�B�d�R���A���M1�9#� u���Jů��#����G�E�>��F,[Eiu�;�'<�&����YY;W��{���G=t�� .��i��m]��Y�����p��\�Iͨ����<&����\98�Cû�t��o��?Uˍ��D�_��I��5�[�ˆ�\�'V��f�Wy���^x��*ѥ�\.�>��n�g���?�nW�٪rj�e�
]1��8W��db�������xh,���I�:�����a>v�Qum�g���֭z�xŃ�YF=�t�XN��q23E�'�@O�>�,�;WZמ,��2�U^[��;^-�wѕ9�IC{Z��s�<��7/�F�hZ{�ܵ�α��rV���|��)�,�8Ɨ��h�����7��C�a��;�=�OC��G���c�P�2�^��c�'=�t�D�1K�������G��F��'�I���]��2�è;��u�.LZ>C��2j��-��夞&��ԛ~;��g��G����5M(3a׸Zb���5cE�]DM���j���W��3� ��M��r����e�A䰾�����ϩy���4�|�X�%�t�ה���;y��qjk�(��݅�1} �f�9������X>��B�q9�pj�5�#��օ�>A䣘NN�xZ�q�On�213�Z�f���[%u���,�Rf]�koˣ_	҉q;��� ��x��}򐁔u!ag������4�o��8؝��~�D�D�\��f��'53�
(Ԣ�\	��hP+�/�K����H���Lq��������$q+�O�/�����Rɩ���,N ���@���~ְ����j�$��U�Ðg6Gs�z��4�8N�^�w ,����*���OҬm��4�O���	m��ak�����uo���$�HE'��b���YA��-��J)�+U��s*��^1��>�p�jHM������x{x?֙��m�Km1I<�/(1ۗ�*�)�)y}���sE��ϫiG��)��"#A��K�#����0a<;���&!p�-��S_�;B%��8t���FX�6zRܴ`A��ڿ.�H�Ċ��*1G�DW����*yf�-��u��/�i��������L{]�>M늽�{J!{'P��ZF��o����K�b�s[Dr 2O}B��֦�� _����1eC;M��C�</�0��G��O1$���KF�
��W��I�R�	���V��5��f/�pǧ�ګ���SR�!{��Dq�4\WI. ���ʖm� Y�3��]�v=Dk��cQL� �f��erroR��k�ck�ƫ�_�#�?R��j)��pq)`47-���xt����Et���)",�`Kɰ_c�pA�Q���'f1�a�9
�a� ���\6"��F Sޡ(:���E\��R�nڹ� �e���X��v�J���	ME�G �2�~�W���&)����-#��y��|�� |�[ͱ%��gݕ�
H�8��b��+����j�����]��V����
_0#z�B�f�?��J��v��'�&&���F8]$!���T+Z���4&ؚ���:Tc�����U��ŧ��f�|����y�d��B�p!:���1�ƭ�zU�\x@ե7q���2L�H��3�-�:=0a>GN��j��(w.��*'�b�	H<D�V�UU��;� ���9�4N-�rW>�t)Y��j��W�ɞ^ZΕ�}V�\*�_�8�Ktmt<X�"L >���y���_����
�wv9���~�9�P�M���A�6�B����z@X�����\��0��XN\�T�����b^#�- ��a�Qo/Ge�[�h�P��!��ۧ������g����uޕW�^e(w��;�ßD���;Tg!w��_�����6sr���Q��^�}�px��gc{y��S�hU�֒��j������
k�g+ˎ_�ij�oc�����V�`:%�5>�&k�.6(D6#h�����6�ܡ�ݙLo�D�Q�J2'�Q����|�yFG�����D4�B��	g��2$r������ ��+<?
��=�U'QÔ����Y����?G)�FO���t9�F���4D�x~�[V}�oƟ=&e�Z%�t�C�3#�Y��	�5�G����j��!@pL�ĥ��MH����"JuK�UH�*�Rߡ��(w����|UR1<��)AYs���,s*������Ę�:���@H3P��h��R
�=�l�;�kJ��D����O�����&�A@;r�y\�s�&�%̘��芁�=���Q8,ud����"5��ˢ҃����v��pdB�R�r���H��V3jY�T�eG�O��[{����6�]�($$�<	ZQ|4
���L���yg��F�8�'���N��Ѯ��8�䶪z��|r%�R�'0�.)�?�3�*��f�FZ��t�ޗ�L �^K�IS=YzǸ���Ȑ��*4>c�����A��WLL:���r�F��Sj� ֞\\ܮCH����g(</%��I��M	Z!({����ݞ�G��e����Rnpi\Ruܥ���A�C��P�"S����<n5U�6d*�Ӹ���7Ұ� ��(E��x�o�������V�������|�L��i5����߸tȄ�0����^��י��!�SMW
�{PNC���x������Y�^�I�m�!ۇ��']�nU��2L���пB��o�KX��\�En~e�{�<�����wO��@HkuxR�i"��]pH1�v��sO/* ԅl���6 �H,�K{�4w��h��}��D�:!���5<�p�p;"�o�������2E��N|�[Y���)�$������|;�B�WlzAky`>�^�(V!�dQ�V-�� ���9�VL����,ְg���l(^F_O�^�~��V������=Nڑ���Ivro�ڥ�e,n�O����>, ,�X�~;;%�D��w_eZ�'H+�jy�&����Z�8䘱������p��A�j�����Լ�7�ˬZC��荄�@}GBq/.��:��q���� ��A3a��)T��G<��{,$���s���0�%x������n��Dti�T�A3w��+/ƛ�g�΍t�6���Pn�{�Ⲫ#X�@c1��xz�̬���a��ql����F-҉�/�>Z��pbǝ�I�z'�X ���;v��\$�P�S�^�'��Lӗ<�,���c�[�S`���
U���x��1��ʓ��=)<������Ճ۽�u���uy�AOӋ'��y�k|�@]�3��,��j�ߏ��
�����ď�����mr�&p�*{ռ2�E¡)���v�pU� ���p�vl�������䘁���כ< z����Cwc�'U�c��A��!a����[=i���!�`�b��@�u�Ԡ!�H}A��.������E��ݴn�>y!��E_|\�a@v���
m���
.ތQ�n&�&��ӻы_��|��Z���!��qb��^�!�N��U���1]#����%�96l��s����[���CT]C���
:�I�,s�5���(M��W��>��v�B���ҕ_()՜g�{6d�"��ۃD�F�	��Y�h�Ғ5J^�s�����1���48�?�����3l])8��H�͚Яʳ�໣�w��Ђ���R�2��8�˼�0A�z�c`������u%�A�bN�bQ��-��Z��]�u�S8���|��&�����=M���x�� �Hw��~D	�d��Zɇ�Nd�]<��h�'F^��p�@�:����V����D��}U�r��k�\�Z�k���q�^��w��u��<oo�z�MԽ��2��&3��gE��W�E̃���ᦴ�GV��x�I��	#Q�]�8�7鳘��[m�$�^���ɀ�����H$�
K 5Ό�	W�y�]�<��^z�A�g�n��}�]*����W�S_��gq͈�尣rW�٫z3��t�	5ִ���V�`�z�~�/FE}d�������׳l�l�W��4>H�v<����U�
� �`�pR:�s@���������@4_RE�,2��=;��,*�t��1�A�GSo5���mu�9�x�W�%줍��m�.
ߛ=!����L�SbN|ş0��j���ΌB�dX��]2��wM���'X�-����rC|l��������{v½�Tn�au꧒n�N��9&�{���&Ю���-�����Z13��n$���9TB��lj�#>T���$�2��v]�{���K���J4�	tl[�r�ζ�,IZE&����4F�}��W}�l2�b���DY�B/�:�0K�tQh�én8�1޴��I�¦�5[)���e	^ɂV�i�-��1�BJ���!W�������9��nT!��9N�]����=_(��e������c&���=�~��yN�k��s�{A���� � <�A��~����MuwP�^���6+�76�=� ���˞����0h�&4��nߙQ��|��?�Ukbrt�yN����AM��T�����*�Ҧ���=M��=�*�#*L2ޑ�Yk��������3���ބ�ۡu�Wj˳g�Ƣ%ܖ_��y5��o�T�g�*biY$���6�ƈ�����XY:�2dP��P`�Y�0NW���K�trD$�/�94[�5��ґ23��}��t8!U㈼p��S)gøMs�v�|l>;�:wn;�X*wa��M�&s_�(k�^EU�H�wH����2i��V���U2Q�>A��Z�&�|�S��$�����C��uA��4�ϙ�L�B�<�bz����Y�0n/?[�p���<�񶵨F���l�ĉʢn�%�iry$采����L;^}2�
'��\��9t߿�ޖ�	u�|YI������-%n��"-�x!P<*Kz�c�ơ=���t*�w�(��r���Z�O�r�^�Vj2"d��(a��f7<؀"�*��g��	������&�+�`�m�qm3�P�,�gD�Ue8'�@��"��P�A�O��]�o����끊˚dED�D4�Y��L]��^;��Z��fP3��xI��c+��in�>j)7�GBB�=¥�ưr Ӂ�.+�z��[~�-��C�B�2��-�y�����q�4a8�(/sz�_.&���8�f�����9�2�ؖ^q��z���O!�XOʊ�_Z�@���'��_�V���y1B63�C�V����ZS��N�i5�b�n({����^�>�Mi���S�>��[��=�c`Vj�or;J:�{1m�ߞ�p��3嶃K`fdq�<��Xn_��f���z�*��JY������P��1$J���S5F�%D����~	=d��HgX�+Y�5�ד���}(���ƄrNor���X�fB�:,�u���TPRjEoeIA��9��O��t��,��G�Tz@&�V����[�-x��~���:���imWg��/�J&7�MG�	�.�p�s�ۺ�ezl>#U�≀
v���
�M1u=����\�\����n;,��s�c����@���#r"�A֮��<<�E����1��{��oT����~n�"eÂ�ʂ�L]�V}�A������ �<2(�����z�#��Wws��5"NПTpi �;�!�c�{��1Esʉ��K��AϜ��%����=��T��;,��]UJ�@#!!�	����<B�P����T[ԛ,���]�)���^ %������]�����$O��\F�,���ܱl� z�!�����=��5Κ&&p��,��є� ꅋ��.��%A�=��e$�Hhe�����F��])[7��Io�H8g���I�0 {��I�S�J�n#6y>�q�6'��'髯W>�����E!a�+��!ه���-*^�BZL6bo�&a>aahi�U[�bf�x>�� X'��h�M펎i���Sp/z��B\	�J�d
��H:7+r9�u�쌌x�$aj�c&$Vr���c�\B�¦��o.�����ߎ�Q�K�h�5���V���{��vl�Olޱ����!�p?�i�{d*�'T�M���~��ػ/f�!ҡ���'�������Yc�M!�.(Պg���0;mI'�C�9��[�oh�BS��]E=T3j�&z9�XI�Wg�j����7�]`����z�I%Ͻɇ��K�p�Ph�=sE���d�0dx�ѱs�zҶ�/�`/2-�|����`G�$�
U��7���p��x��\���=eKqg�/�/ё�2���5����I=u �蛩���^$A-��Х�v�ZJ�?�ɬ�*V�B�_����o������;v�z-�h���$�e�\m,�?<0� �w�;���P_�	=/�<\a?č���U0��h�w�>Zs��,�9/;�� ��.�p���QAƆ��~��"�V���5̴�b����!� pR8�O�&H�`�5-!wʆ���W#��'�J�!p��r�C\��&du�<ZJm}�W3�c��AQw�Y�Z��X������'��W;�_����	�cŪjHc�!`�2���v_�C��R�e�_x��2�Ңl^	�@�����\��c�n�o _&G*��嗉���2J��ʀk��!wS�F���`��\w�!�ŀ�ymO�������4�硞�eEmC��z&8D�ƫ8� �Mid��I��v{Z�:��Ož�;��X���^蕶�Rf6�W�:�{�>,2��w��>U��&����J��)�j!���Ѯ�ч���$�P�?b�[�N�D���>�ع$��e�6���W`�\�}�%d���?ɫfܕ@o%f%�x���_ԃ]�s��k}��aC&e�����DAw"��݀&>e5>��|�,��-x��h@�҇i����CG�9!E�HV�d-�ߦa@�+_H=R��G	�N�y�Ł�o�+���81}���a�#C��΍H ìζ��' �5�J���A�bX�Z�TŞ\T����������qc������]��d�X�Oa"��84LH|�sr"��ܯ}1�yM)�8T3_B�S�c>K�_k��3�<V�!nҥ�_?�k�LԷ�О��97x�H��N��Y'NM�e�|�ze�0�aF~IV��R���s�?5�s>Wn�i,[�+���+�*]C��޼�v�Yg]8��&O�]��e���{���`{O��:�x �)�@?X��,I���f[��b(v���a�ϯ=t�Ͼ����;��4�4�mG��l��G�M�&8������._B��b"d�u�LЩAW��v}+ѻ��W�F�po[���D,z��v[��q@Q|������s�e�aN�Z���G��Y>(�����Ц��P��
��?KN������D��rₑ��5��4�p%n"=�n):9�p6<Yi�|�!mO�O�Y�#��沧>/��%�) �`s ���Z����j0-"8��H.W�z�C'���mT6٣j&�W^m�B��,+�z��G
�/�w����X�W�B%e��n���`a<�Ŗ��ZX�y=!�p�rc�]! F�N�kU�Upw[��vL嘇�6e��.m�[���K>e��������Ƶ�E�Ϭ"�,��ʋ�\d~E[+-��<�+j�:W�4� ���}-��y������*^��ġ��2���A���,�:/�����eJ8$�R{�%B����X*�.�a F���:[�����c�Y� ���y��]�_�\r�C�oڭv�E�!��v�������0xQ���I�d��(�ҟo0�<˪/Sɣ�!���M�Ԝ����X����k ���_���bLu�6�j�m?>w��ar�X?։b>����'��>��zYɽ��x��w�n� �#���="p}���yˤ��m4��*�6nֻg__@ϳ�U;昻U#�l�$�'����Rȝ��L��Հ|Go2����G#t�/�3��a�=���rf�p�Ғ.5�ռZ@|�͜Xk�j���	n���W�3������/���}|t���:��b1��i��Ѱϥ�R�c���;�uv�7�̋p>N�S�4�l�?��x;w�uh�7Q��\6���;I�q���;�)	/�B�
���z7�5�@b7
�p2�U���Y`ߎy�U��lĉ#�M�@6����+*@���7�?L��D�R�����o�	����z�� "�.��|U�E9�5�G)��KWR�X$�}�%Ŗz.�e�a�$xL��IZy6Ǟ�e��}
��xQ*a��$��-¼¯�nCT�A���d"A�jhZ[gmc4�G2L����W�䮈�<ls���g��s�����<�����k�7)XI���Gg�b�iK����ޗ��}�5&�ð#�娑�y��/�8M+�R$��m>��}`m0?���nQ<���d=���uE1�r��͋2oZ6����M-k@u��&84��h�r��|�k�"C	�D����X/�E1J����j�O8�xn���[��[���X��r������&���_��Y��Ln3=����vw��h�Lc�T��*�~&�ioK�6on�����a	{���p-�9/ü��C���4]sk&jd��WW<��Z��4���-�rAl����v��&��D'������݈�_�e�j�W�O�}J��$	�_�R$�f�p+B�H�I��E��&�jX��'Q��U�W����,t�Z��"託�D� Q���F8�ɑ��;z���dl2���W�5�6��Gl�T�E4��2�ܻ�E����ը�yЈ� HA��@!��0�CD������:�z���	�ZL���eD����6#ӊl�l�������D,�q;�i,eT�5(�)�[�yj���T�ǷS���w�ͭ�tƻ�.���e��&���R��`�q
]d���\�\�ƚNF�>'eo-@.��"��p��/�+it��7���~Ɗ��/�J�K������P)7�����J�$�p�\��weǫV�B���W¸�~&�d�y�Cv2�p۩^��Ȏ��v>|������;z��r���Ef�-�a�t�t�[�|����b�@���4�@E���:q�,Ze7>���LP+�$U���t<'/�nKu7�T�P�B�1� ���;E�U�����Z���:�NJ���
E�f��]a�FA]�� �Fv?u?m�U�m��<��@�}�o�r�x~�y$\��q��[���,R'�h���3:J�O����+�� m�]g����8,B_�fQl�ǉ �^ޔn�X:I��w��'r�^�l�J��ָ? �6��Z�ᶣ`�`��V*�*ӟ�I;4���N��܈Cz��/��C��Ud7yD}i�L�#T��7$Q$�Q*'�2'����]�����g^�&��	�LD~�M�uD�y\�}�V��h%�O���-���{1��ub�7jiٺBķ&kfvU��T��F+&���¼�9�Q�!��gǾ��s�}��b4�m�ڞ+Z;����'~�D��'-$a�C���~�h�w��g{���iO�U�����n��
�1�� \ͤtd�,�/_
]:c�R�9�lCI�
��S�]>��P��	�4��Ő�B�B�s �H��$�GxB�@BՠoLm�����r�+�m�Yz8��͙�dr��;��OXc'Y�X$�ȕ����I�h8Z��#y ��u��߇�)n9.he=�MG��ڿ�����FQ���N���
>�z���b��1_MXh1�wb��*Ҁ���v�dnm\�Tt�g�����3 "L�TۭQ��o|H��'2\G��Я�).7\���.�(g�j�F
�]y�������Oc���9���L��;v@��S�#�X���Cb���$G�=�5%9��b��k,�5�&��=�?�T�OP�����b�����2��id��(��r���F8������	��2S�y�Xq�e��G%�:�A<��:M:.�����Y'tRW��] ��7T.��q�R���G,�pG��X���N�q;��e����J�-�����K�f�_�7�������C_�	՚����I��a�Xh#>�A�l\I�H����r��sz�2�1Z�l�#�&��zh��r}����ip�����)-����f���ז:~�H�3��% R���D�^U@?�76]��	V`�I���ֈ�Z�&*H��W����9��Q�q��|0����2D�#�fn�j�4��r�P���0;��3/�EUH������{��LDW���S4 ���Zr��x�`�u@aC��%�u#�p̐�`'��_u�1o�Y1��w�<H�Fz'H~X����qM�5"�l�(-�MKA�#R����>B]0���>��{��ݙaQ�U	�ò0������/�5����\NQ5���3�)W�X�^2���cR,��$lMAQݾ5���PSL��=�
��? �҇K@��/7Y�50e�c*�~�_��{B|Y�5§ۡ��ё�7]�+���R��ǣ��}���ZLٽ��>W~&�̞�\I���8��QT�,6�ck^Ѕ^�=�K�r^i'<��ܝ��Oj��:p�h��J�h���%���!>�����a[�< �Y�X�/�����9��hS��* �	���2�U��1�]_��tUo]'��(R��J!-� zP�,9Y�ǖ*��S��!�̺�%��s�>A��4	3�v|����/}�\�Ӟ�hŃ{����Q+F$E�bh ��W��o�'
��Gս�s��jS�^�#��Iv�����C�J��>+�{8�`�3���/�+侧YD�j$�~\�w��h�
-gfG��}�՟0Ʊ��9&� �(k,�ݙ���y+(	�Ř]�>�5T���3h;[6���4����3�tB
GQ&
�R}GUG�Y���g'��:�G�
�������v�q��8��E�o��Er�V[�	5����Q�:Z�^'{K�L3劏��i�{G��@�#�k�y��`�Bw�;D7�?����xH��Q�;M�sOS�EC����b�H.
м)�|V�ք�s�'�s\���7	1���F�/O��8P�R1'���STGl�!�R	�`�����.��J��sJ,q���o�tD��!{sI��זi2���{�g7���:�J�r�}I�P�AbCB��?�^�~����y?�E�㿟)P��^�4���#p*�(�w�NZI��e�b��c����� onO\Y�+�P}������æ��������[ӝ�#=U����*r���f���4��.fo��E��ρ�i�61�+�7�����s4������.��1��Wh��k����aӋ@�t�0�T�%�H����--I�8����mJ��b�����\����f�ޤ;��]�e�9M(
�0 �79�F7q�Ԙ�u ���+1����d`2�����`�B�0����qF��L�<�vA�a��);�.��F�Ӵ�@�2�'�!�{~���� �K�5���u V���v�.��U,@��wQD�ttx��[�q��t���$�G�8���a���b�d��?��|H8�Szi#�� �p��T4ƀ�u�]��3z6p��Ò�T��L�k�Aē��f����Yz?܋3�t��Z,чL%�4g/[E�CV ��zl��0|�@>���( �uпojs�#_��4�M�4��r��"%���2���4UD(A[ά��7���a�J��H�c�\������`Tb��jxd�Q��\��2V��+��\��
�cRL�1�30]�R?bm	
����W�o���H�J� ��Y���<������}��A�Ϥ�\a�Y��	��������uP�R�}�o�9? n(���Ϡ�kK[J=�G��9�^��F�c R�e�;� ��?{�T�A�bm-S�mZfA�T� U�� $4��S��}AI�*1��k�D�ub88r���,��ܯZ链���6���� J����N��0%+��KQ���ڨZj+$�6�a��GQ@[�U-y��qfz�����Ǫ����L��f�����W��m)����Cq=���w5�����B�b�D ޿����eQvn�Rv^un��x՜:�M�$�=ג�B��>�A<'�q`C��#�cQUK�vϽ�묱z�%�'�g��w�T3�gՁ����2�� ���Ä��W�@�e϶��TZ�!@SJ�dF���$M&0i ��ݛS���Ô�������^�<�xA�3HK"���P��$譭�'�I��ܯL?�Pug�|w�0ո3�t�ݼ�Ǯ�;��uf�t뱪s��unw~bíQsG�����#����f��}6]!۷H�`��д�.E����#��ѩ�p�Y�B<����'��9d���\�\2o�:�ۋ���a�?��)&:�vH���/��6`"�%j�~[�o/�ܞ�h�v^�c
�b�!˅�PfK4��2tl
8�����:	'�lx
g/��~��!��]�W���>  %�A��ǇYZfvU��'і�k��Q��Nj�́6۶�ϒ�YG��WV=�;���f�>c�<����S=&��r*��"��/�|M2�@	�kڿ�n�d��F-����XP��`)FMu�Q�$�r*��� >&�͜-b���4�נ�NP��/���@GZa4��A��:�$���@���ߊ�{Jc݄���s��e|�0�˗^ſ�E��c��'�V�;n*�^z���������	�j��6���v��pxՒ��h-F]����'2��Q�qsgM�Sh�e�m��R"�E�M�(܃(p�ٖ��X�<�&~oR��F�b�4�6_���2Gܽ΄��4��F6��dׂ:g�E��i�ަ�H[(b��l@� �#��%��R%�SQ�FM�&4�]�_��Ӗ$tܤ��7D������E���qISj:ف�	M	�3�,���a�C��N�U+�E��6�\���B�)>�	g�>�t�-]v�ק�ܟ�b؆�=�7n�R�˻�	�l�+�RN���5����b��/a	���)��m��K��J\Ͳ��1�����I|Jʉ��y��ʰ\�1����&+��6g\�F�9֓2T��k��Al�ѯc�5l�l�?(C�%�R_MT0h�w�r���i^U졍��i�J��M�N���8�'}8��Q�jC-��<|�L
�C0j�;��&�Gn~�.i9�s$�sFFdT�;��F��ZNfzdw��Pb)3� ���I�A#��;'��jd�&��0-2��G�{G;ǛmVZ6)z�q`�ԑ��`e�A)�����?�T�~�ˁ�%c��O��ȓ�r�Y��s[)�;�L����Ҡ����,k~X��/�+Q�m�?�F�\孵$Ow?��odWO����y�n"�5B�ݧ�;����~���Mﮅ����XL���9]��F\Bu�)���+7!U\Ｈ5�u��/gT��۟[��W�&�+�2;�pԖI���]�% ���v!ɴN���S[�jP����`_�L�\��x<�+��҆f��丢��A��j=���#�Jq���M4њ�| ��%GB9��"�!�z��H<��8��-��n���E���۲��U��^[�X
¢�v�5F����!�G)����#%k�;pH;��iQ�H��=� ��W�O�p364��L�)���E���;EH~i���7��ML,�c�j*^Wj
����7c�$"M����LIŮLrÏ�����W����bj+�+��Rd��@� ���ӯ�&��N"���hS��HK�'6�,:E�z��'�l!���u�ν��
�[�6K�]�:���t������7�1�HcWMDu��m�d�wћ���v�2�5\D�R��nŻ�lhΉ��VY�'CL��Ew<�a��4�RK��l��	Z�f&%8�����E�齦7���U���1�|�{`Q[fh��]RA�spm �,�XХ�՝5p*�hH��yA��'n��~w	�}�O��#I��Ǒ͖�'�s��xaLpP�'�1�q-@��zx?�.e]&SC�	�l��n�.�]�t=��p���]@+du�'*=���YTV#��朗�g�U����Ow���`^�9a�n��^7�[U����>�R����������$�̄���(�v�^��Jڠ��V�c�ð����|���f�`���8C����Pl��d�^��s�c�2;�j��YT��z�5칄ذ<�)�3�zx�|FQ�@�l Ҙ��pym��*�1�rD&Z�f��}0�昫)>S^yZ�^S��P�۲D�{5�zr\���'�9� �����F��]��8u���eJ��S�/ �}����fX��O2K"+�5MN��G���*�2\�Te���k2�+zsK�����a�M�W�z�c�CA.�
W�(1�o�.ہ�z�K+Oz��3�A_!�tJ�[�����4��]�ΝR
�T����c���?�H$��du��"�P��x��t@&�+^�@0Z���쎚�j#�^��x��g�7!�� �Ȋ^�Ha���o�.���rݠ>z�]�J-7IT�h��Ѻ�De�������E⬐��`��l�ٍ�����aYV�6������T�S�߲t��6UC)ШN�v_�΂~W��CkGY+��XX�'��ş�H���r�cH���kW�2�� -��i�vOs��D�������{�A��x�D���J���Di�vy��e���Ċ�\�/19ɨ'2��a+B�e3,�A:D�&�*fr�4�����)P���68ӧ4�����Sru���e�Z\o���W&�a)$*p˥��%-�ă�˖�&��.���J~�у��������1�\���;��0}�9|j>��VB6갴+�g�3 p����h�G����Q���W�=�6��泟^.�j���1�Y��|dD_6yq&b���u�@���q������c�G"�&�,�̮ӚN��.�se���{t0꤈:+�p�G��I��F�jϒOsCsy�[gp0��m���L���qiT�]I��\�#��AÆV5��_"���q,�9��tۡ��_Z�����7p�v)g7��~>7?�8z�5�M�|�?Ϋ�-{�B׶=D[�O~  ��y��D@�CR�J��Bd��J�SȅJ�^��$���@��m���4o턼���r�7����nJWFο2�$E�Vv���$^��&��?���t�"\#��;��矚 ���F�
���x�~�	k&�*�4��t<����{�\�A�p�3�b@�??��ϒ�f�%U�٪{8�L6ᇇWSM�EO�/�b`}�x�"U�B*^��G��s�0l�ں��gF5�LY�䝒��$n�]>�۴�q!���ǋ(8�Go20�e@tq��T�n�fM��	�ypB,�������b�4+m�d�9z��5_�q��vc��JZ�f����2�Ӄ�E`���Gu-۩��wl$g�_I�d���<�ԧ���N};g!9x��?�|��.- F��Y�03IO�A�vu�nW�"�[���,p.OWѬ�(qy�jK���0Tc����� %u�c��[��r0���8G�b�$䈚6I�s�9c���	.�]���9M� ��4Ypj+��UӤ,8�_/g�r���c>��U�����CtSz LO�S	eo�I.�&�(��2�,Z�M�`��n�to����������Ս�gϷ_`�b8��e��,4���8�W���\?�gˬ�^��)��+
Z�J�����b!:�kL9&�Ü�h2� H���ah����f�0��X�ֆ�/\�΢nmߎB+2�i�y|R��%�Ȋ�}JgfV@�3nI�k�D/6��6'>�����P�fm��7��C�*k(r�������b�r��\Xw�����Ưl<�.�B�4pK��@�1�܉6��J�����Y�ڃgI���U��ɓC�E��CeY�U��$fA�1�h�HI����,J;�u�$&�8���_�� ��C���3�t������V`Zc�����*����*?��ւ�i�+r�D�'R���>����j+�I<`�����r;Q�/�����k��Uu+�5mv��l �Q@���n?��ѳ�g~ƾ:��>(����9SK��U���<G�7���
��pa� D�s�%_��������٩�*ť�F����Z�����yI�q��O&��\}��UE�Dg�-:*F1�>i�d$~,jNJ�V�#��e�b䠇��ф�Ⱥ�@!a�H
�=�oi���i\(���է5����ՇIl�P��I~����{��5�y/�͌gf��Xݧ�_i�T��f#��9C���1]�x��
���ӆ� t�1��R�7������"�k���;b�$�ZW��P�zQ���@z�D�{;���aY=>#@�ms/T+��~X��â�W����ڬw��l�;�!��W��LP0Cbb&]ԡ� ��]wsk�}d���N'��E�7�䯵3*�b*��>m�8Ʃ�(
�@�Q���i���O�/��|�w8�F[��e�<[��%O�ڍsd��j�љL�lp�wZAU3vq�����{ֱ�\��5>5�g��Q"!�5"]��:(P� �t�/�%�[�a�vs���nbr���t�d��1}@�9D!���U3����$�E"�.�_�<�ffa�� �*��[{���o�w{J�J�~��Kei���س�����=,���v��=��i�=H�9������[���������.�eF)�ˏ�ƴ���<�ZNO˂��v�q~�c^�%k՚���E)�oʏ5�;��שH����dl�O5�G��#��"�v�6�ma0�O@��wE�臙��A磱�`>��a��GF䮬+b4��#�f&nŨ��C��x!P�UK`pĢ�'�Vp���L6����Z��E��_�5tz9�r݅���'���<9k �Q)tl�W�W�PV�r�j��-�K�)���	�+��kQv-�����S9���N�U�J��ER1�`�6��4��G*�TIGG����bY�]q
����呟�os��!�~~��G0��	[��4�,��$Gj2�`�4�u>�n�U�)b�,n�,z����Q�u�D`J�[��\Ϋ��B.����|�+k*B=��рa(��g�&c0�O��@��g|N{(�-~4���ķ3��@iZ��:�1�όɀ�a�Z�4�A3��e��{���:Ӊ�g�phOt)�4��A*?�>�t��D��7�aZx�����s��y�� p'��>�9������>'��E"�&j}G�u�:؉PzP����J�X���u�d�܍:�}�K�����<DF�]�L���bW��Iz��E&��5!��=��L�1 FɅ�E�OW�q�0)�;~��L{�I-��;&���i�"1h�|��+9�c-A�������;8��R&qE��_�7$��~����Rs��/�*����A GsP�P���HkH�SA������]]9�k�u���a�Q&9X�{��p�j�<5�A��䀻��u�B�#�o�̕��Q?���8�N:̃"
��佌a(�_�qm�[͟�"��uu��b�{�&%,t����5!�6�����
�Dy.lgϞ��V�G�"d���r�����L1'��ΐ�_!�Qa��� Z}�q��D�����"�~�bN�3�ĩ֒���O�Dh��!I��:���uY}��O��X(�]sZ�yP�>m�/�;Ds�o��EЂE���-�}{/����<]��J�� s	{F������o��0��u��a��Ϥe��QD���U��h�D��٩ְ3P�e�i�S�"��	�������"��v��G> �=�`C���f@�D��r-˶]kŹاӭ�R����U*e����gM�W%B�8��o
���-TX��_ ��5�V�i5^N�0��)��J�umO�+|�~���U���]��jD�_@>���N����%�,��^#V�w��A��'A�?a�x$�F^B��o4JՀ�N�c�?L��ײ�Zy�\�tx�曄!�H�!�uh�˚��A��Ӯ��4y�"])����l�W`�*��s�>̚�9�m�N��5���g_C�!���\ëdx<NL�m�U�C��i����A�L�K"�H�����k�$���n&���Hw��2����Ml�f}�T�7s����PD��}Я�Ϡi	Bբ)_�M����q}��#��{A��l�-�����V~EY$����eu�?����Sw$�#���K��X\;6�3�5dSh[���ji�p�ݹ2��u	c�W� ��ƻ#����ފ�R�f\o(}YX��\��.]�iMû[9��(;OF��o�֝Q'�ǲ:����o�2��E�L�K�N
k������Pḿ�P��������_���o�ޠ}�V�0Tb���i�f������&��*�('�����&�V���Ζ8/R��NP�7ӻ7���k6Cɸ寡����g��A+����08[b+�w�"���0B�
H��u�LM���a�����-��bQj��:4����;K����4.�S_� ������l_'g�E�K|�j�˳�n�2��P�(o�+���ޝdC�C�7�?ɠScz;G$�⇝�F�cH�c�q�-Qh@%����kDW�������0�7���-���ּ����Ç��\�(��� &W.���"�?ގn��H+���?r"��-R�_�p��y�z,Ƚ��/c�W�|�?����Utn��H�P>��vZ�yOt�}y��&���!�'Wa�����ir9�,�^����	.D��$�W��eTe�j�͓��bn8�M,Y��|%�����E���{����)�5�㯑���b E���������޾	�fI�S��d���5���{̬�a�=���دUV{=��Y�?&Rc�	���*>�����cO�L�s�Qv�&�/�=��RS'�|_Z��j׵����c��;ơq"`J��"ْ�����3���[��y�EFYu^֍��Q�����>����/�����]�r�[�E�����9�����r�����]�%��r��23�t@�B"HL�3����2�;���PK�Y��:�צE�m�|��Ő�����n���8Z�U��n���9���B~�h������K�1D�T/Vǵ��td��X?���u�ˮ���+ѣusm�1�t9\ȹ�CϛV�����k�=�H3|�G	�JƐ>�&k�����_����%�[��ZQN|�-��#(� ���h2.���C�U�>۪p‹�
B����[1s�*�Ҕ��g�]�#aD��K�VF[|�sy��=�*����Ol݃	1��S��D�3��e���ڎ�}"ͽ /=Wcr�}i��_i�L_D"�t�~�F�Ǻ�l��ܟR\쨼��+=D�z����A�~i샗WHS�j�fPp���:5���*���4L�=��/C�i�}�$tur��g�S�+{��	��K���hU�y��,��B�&��:�d�;a_���6ays�ED���o��;m���h��^�K�:Q�Xʝp�����c�Y�tK?�ى��_��Y>�SwL��vY�Cȗ"͙��9\r0�#�bp���CB��&�����	��X���K<�Ĺ�%~�*�K�.I�t���C�n���)R�rr��6�V�u���8����.3P}\��Õ��EXfx �W���)��G���d�U�{Ќ%���$�7Q��4OU�پp��ɑJR?H��m����b��rj+�Yh��aUq���G	�?UR|j�V׊`�^���4��m'�F]�:c<o�������~W������5�oVf��9��ۭ�P��lJ������W|A����8l):�I���M �V{A��k#���x}�q���L/���'P����L�t�R�>{q.N�䆘���T�O��3�4��I@�G����h������K����t�8y�¼z|;e;#?�k�+����DcV(:�|���c&o+*�co�mi��-����^��)r2<��5 �份�a"l��>�
��Mx�=���<� ��VP(�ۧ*	�Q�p�c�64p�mU�Y����d��Y������v�����ő�~<���A�]!��6�h����dZ\��[C:\��a��n16��3-�S��&�M#�����L����NB����Ά��G.��s����M:#ئ�(A��	��h��H*���8�n	��Ve�c�~|�4ɐ1�ZEޠǫH�1[�&_c�U6m�Y�f���Mq�C���2I�Ԕ�`2�����g����l�Z�L������M*��lu��Z/=^�vC>��nS5{�)���
'E7�̷��֢guoX���>u��?��A�N�.���==h,ǐ�Mu3\�������D��*�`x����b��	�H�O|�
��u�fXZ�0��� [���zn�!l�W�8
�c��d��b��^����X)-�8�Q�a���vd�k�p]e��ցL������0␘I���h'��Ȣ�>�q>/Xx>��� XCoI��o���|�g�����g������mMH`t��[�O��6��\� >��UG�2e����N��W�nChՔ"q�6��]TT������S]&��_�1�U��H�9q�E$QlGfA[&���&��@s1+1E���K����e����ʱ4�E�e�	�T�ڋ���a�:m��i����k�����z���<_�vǅ�g�D�d���7�-����DϞ�ߎ�ոLbI���蚯	�8����=n幹.}�Q���$��1?!�����n�����^1K5;������� �?�\@}Se�>�cRp!6u>��M��;\>z�������qw��>.p��Q��J8�֎��U�T�wGht#��?')��2����A�z
�*��,�+����
HF�H��k�!yK7�4���;1�f��4��O����~��]H�����`�FDU�h��?��1�
��7��>bW��20  ��T�9���S:�:�¸\��)/;�ά
|��!�+i��g����F�o�@���?
�3N���%���O���א�����-���ev���Lk<�ɥC;�(�P�k׭4�$�5�>�[�?�2��˖N�Ʃ����
�	���h@" yZ�L_�W�ĖW��J{�����W�������X�Lܩ�����ck#��`�ԭ]bl&1o*]p�����tL�X=2�h\��m�fZv�[E�gOX�sF-WgB)a~�d�G��v��>I��gxpA��3���j8ZM���oH5�Y�3��ś�b�N;C�� В�T e�Ol�6��C��д=�t��\e���_uu(�~��W�z|q�j�h�?
+BC)��hR�B,�c�b�Z�4�]�Nm*�KoR�zT�vM[�Ly:_�8Y�@.f�y�2F�1-��4h�.+̷�u*�z��
�C���
WxR�{��H��g�Eq*Ĕ;�I��瓹UKs���`�"�Ri%+�_���"��6 ��Sa+7�|U,�a�̼��L]A8R;s�ı/�h,�<�$���e6t���6x�B�)%VӁ�w�����2Ȋ����8�=8D���.;�h�L:����lqūv���.^G�k�!H��؋��̹����[�����ל�'�x���J���j�i��vD�Ƽ�y�2���!9���C���(��d��� �����m�}uLFu�ntwQ���(�F��\�}L\����<�'(C�a��.g<KL/��5yq�@�[��X�ߢV;�:����!TC�f(�N[��?M��6�8+F�}X��G�w]:����t��2�t�{`�I��������ga*XN�#�ꣶ��q�H6�Stw�s�k��'V-t)G@;;�E8�uZN�2,�YV�eA�.KF�!���X_��G��_��JwȬ���5��J�U$S�2��W��/r3���l��7o�;#��_R_s�R���xbk���g������s�{z�}#����L�}!:��~�]
,��h�T���)��X��4}4�ˈ�.�����]������=�8��t�C�PJ�b;���;���������!�v@� <Y?��rf$��)��yrEr��Np8ɤ�����e�^�8T��,��]�t;~�.��o��?�gz;�L���'n6�ow1�h �3�W(|8bp�Z`H����V�ml��g?�m^Q�(��a>G,[|�Cs��A��~�'ybϙa)~�Z��ɯ�9z���6�'��ˎ�\9,u��J	C�<��b���q�T&M̘��5�f�>���D��:�9��_HO[����C��gh
 i2'2s�mղ��s��	�]���A����i�aG2��@�8.a��Z^5�oMܯ�9疲w��i Br���͞_	�^5����q�>�q6�{�h���T�\"�ɵ$�?�*CHf�E���e�}�-��Fl�hA����ǃ?�A�:s�%�o>Z���t8�,�7�6m��{DQ"fu���>��+��`E|\��촡�j��&�x�[�Q���9&6mf���B^J��\�+�\N~����mف�Q�G��:[�н�&�2#�����ʃ��z�W�>�g������f݀_1��M�/ƼΫG�����b�M��3>-H�! Ng�1�S�q����h'��*l�vƞ���L��[C��εYN�Βd��fF������p|V����=W�����;+ג����*�/�q���Ҙ��iv�W���Z<�"{�q,1y�m!O�Vb�/��?�.����ktbV�L@�o�sW�N����]��p)Y��u�yZ��R��QR�IrB�%og���p�6����9��n ��ފK��x'�?��2'\��c���W�%&m�v� b���u/y���S���eY�����Cv��L��=��4�1y\��c�.���r�N4�	x%Td7��y�ٸ\0����d���@[9��s:���A��k���6_��ī��jo��Kpv{�,�I�J���Ok���?g�Vg���^V^��ɧ\Ͷ՟1�Ȓ�8A?�� )s(*d��Q��t̤&�^��}������m1�n��ICsC�g�WL3(�����Ν@����U8�� Zi�IF>�e�&ɘb�=����CTEX`HM+RpD�2�T����z飑I�y�˓yt��;�?��p!WdDu���
�,�.��4n�[��W�=�n���.ǟ(F�Õ��1Hi�"��0��9N�@���ne�E�dVxO��aM�6�>����t�+Y�[cA�KX`~�l�Y���c!)�ՙ�}1�N�vT���-��)��~��.-���Pw�+4���Ϗ��`�L�~#�S��L���y_Ix0<-����xXu�xq�LBg���D���B1[[�2�ЍS���4�b��f��P��ri�dI���+mͩF��oi�1e��A�B�TC�$�\�/&�w�����˅�3���]��L�P�SQ�3!���r�cp9��d��I����OR4�9ӆ <{78��'�˱qF_�j>E�i:M 6%"ޔ�/tP�o�D<T����q����?*��r���Z�MƐ�PY9̓�bW*���r����Er��ш��|{	�d����q'�q��AVB�>ʷ��2���������5���i�E��Н���+�)��4>?H��o9�@;lxV�_g�p��n��hl��.I"'Z~j��J�{=~!�S�ލ�]������ls�2fWrE�<�@�H��]]�a~�@�����3_�}RtL���gqc��m�]:��AuPO�J�4lM=��!4���R�c
����E6V�&�������N--�1I��2-�9(�7����J\lloى�����q/�Fć�L0,O̽Z�I���S<��;�����6q
G���X�d0C~���3lHV�4�H�h�j��$s�k=�ڭi�+��������]m*Q�̔����$rV{d��1^S��nwB��Y����,�P��uL��R�7�?`-��յ,KǗmߟ	��iV~kQ�ES�����x�{hM�A��O�&]A���Єwc��κ�_C��<�L�ujN	J�zwZ��C׋���޴T����B�t��H��d���B��Uwf����X��L��>ʲg{�L�o5�����j�5�%=�Ci��q��\�,��g�bd��;����Tsw���R��îĔ�R(b@�S�v�K��ř>L�����Tia �JF�LH2n������f��.3���:��`�j� �S{i��8����̥Z�TQݦh/� _����Gm����12
VJ�L��f&To��0#������_���%:������|-̔������[����j��T��%M��x�ca��'�}\�ރ�9*R=@����@K��F��n-#� c�bz
3��s����Ym��J%z9�ʈ������('��!���E�8���pmo){
k��+���+�#�t�Y�K��=]D���&���52��Q����6��b���g��M���I�w��e�;#G�ʇ���s[zNwvy�JL��"��4�O/�FK�(-t-*]@��K�����"R�_�<"�;��[�ǉG����1W�NP�)Z�p�?u����j�
!�v�z���D�^�R��z�@���G�1��5������ZFit�s�鹏�!�
y����tD�����ﴏ�D�e�sW��eM�z��&�,�愷cYfd��]�������3���/U8tT��I�Y�Aa8�>F\�%��l:y�k�~�7��W�?�/Y��΂_8�.�G��M�)3����px�B���^J�=��\y#N�Sb�m�DB���N�F]r�ͪ
�j�p�YK��.KI�v��Xu-�����o���-%���'�;U���w�k]�Ŧ^���f��R߀�]a���Hp���/�U'0N�e�00e���ެ�%�/���l��7}:���}��9E9.��64;�-�^;���"�璜�Tp�B�,J�	9�F�uo�t+?J��(�Jzf 2����M��?6��BUy{gl1�ځPU ��)�rQ'���G{̟�����)��鶃�d	�'Q��P�yR���~�>��e�l"H��
�i�cK�ݵu'�a���i�I��`���3�����>��0���s���Sc?���i����'��NI�jI�*����Fv�7�j��w��������H�LE��ʲHJ��C����v�f��9}��|Y��s�ik��4�eG~`�7��Df�F�6���?��ڳ��T9���z�s�&_��97 ��D������Ƒ����������D�L���[�\�x�d`wZ�)b��K&���.�ʚ�e�
ǣxh�HL�e�Dx9x�F,�0�M{�,��\��{的#d�|x@Iᖼ{�Y�f�.V��g���ǝ�h5�,
���4��ڜisCH�����+:����+>��  ը�5�M�/b�3���\�r>�*��/"0&�D"Ȝ���|�is '��"�&���{!�ڔ�X��NV4$�8ߩ�d3����'�
�W������e��`����[����iM���n�_~�@+7uL��NƋ����օ:9�����`�Vt�>Bz�jv]�^`����6�B��	T4�b*�Ѩ3D �I�z��?x~J��}�������{c_�Ѡ����h
�+=��k�s���>���-d0��� �H��O#�֓��
h����T�7,��p˕F�K�x���l/<�cQ��5������V&)J[g���C��{M��!C���}ի�٥əzV3ŝ�}��U�K�׺8�����Ym	T���;���9R��l]^W����&!��Q}鉛�(�J��`R���z�ЏDAŷ���
��B�.M�|*u�����
Q���W`�mG�RK2�w{(8���to��6���y��k����8}f����s�րQu��2Aju������*$?��F�g�q��O~z��M��8g�n�&}<F����������6��ݱ��[���3Ӄ*'�)~e�s�Ŏ�}�� ���bK�,��[�\R^�="D�с`p�\����6Z�����KX,�B�~u�� ��G����nëR"�C���Ś��(�}�T��-Vcr����#���'8�ݣ�9�?�19{�����o2;��NUK��T��Ӏ/@�	�N�J��5��<<�|�l�|6h�VM^Ψ���q�A"�v�9���r�8�e��~RٯV���Ho��n�B5t��G����;�b�+�f7r큳R�l@����^�V��=K�,����ř	QAlr{��+4R49�U��w9<��X�o�Ӟ�{T%���a�����af���VQOX�aA�:<m`���9�q�7	�*w�������xt÷��U�dw�S��+�ύ��`i�:��\~Z�Uu��7�pIKZ�IbP���(�5;]}/.�#R�����6���5R�\ڪ�]^}�Xyx�2qA�Uv���Ymd�+{$c)t-W�ò�~P��< ̑��̋JTC�$�<ǽn� �$������%g�!���<���F�vW���ߵ�u�z�:u	{_��f&����u_*�mڏ@���Ck�S�i/C�%R���:v�!>X�= w�#��־�d���g_>�V�I(s)�uŴ�۲"�L��7�4�Z��]��w��j��!�ʠTv��{~�Vp- �`��Z&�@[�v�7���ƒr�3�z��{��ZD�T>��ox8V��-�����`�vBqQ�B��.7�mԈ��12���G�s��1���c��G���P��,R��"���J6��I�lF���|�69Z�_�y��dO�,0�G(�4��(�y��ס�A�>ۘ��K��
Rю�������g��OgKSѮ<�v��L��^0p@���SU�� 7�N�x�oy�o�MG��}e=�g`탙I�nD�8�Yk�W�_� �3h%u{�bY�� 1O�~8��!5te�v�J��2��<\�����;�b۫XR}7����������=�X��ʅ�ߘ/]�C�I4��]���� �}��<m��C��9���S��x�	M9���ή�D�b�RV3F�&��mIll���ކ�-q~b>aں�6�ֻ�@�9d�냨~�����Ƴ7���b����|��<�Ou؛2<)�ͨo|'B^�9��\���^"�B�"��as[*���R���Kΰ/5߮�a�����+H!Vɐ�a�c�Rjqµ��鏣j�"��(��RY� ��:��b�ϵ�;��B���
����%��j�oE ��\	���o��m&���10�p���nc��$F\_�x�����Q>����c�_���Nn�P8L��Մu�����MQ^�
]�o,|� B �e؉Y0[�[c�%�N������ E� 9zF_o	��+��V�Ę��uHbYƳ����<^��u�]Հ�5�H~<���͆�����?^�9ϩit3��
A���������`������}��'�b�ߟXR4B5�n���	�	��+�R���ʠ1�ߣ�q1g%��ҹ����i#�n��ظ!MRU7��J�݄U�j ̰٣\i�)	A5��
���"69�l�Ǣ�m!��O}�G��U	��}��x��U�'�+-2���'dD�0��u잎0+��?���Z�ֺ�&����� 7�=��Z��^�C�|���DHE������C)F���OQ���6iæ�>��Kg�?<*0�ҧʥ�6R�v���үM�J�n��Y� �d
VO����O�Fh�̵M�kQ4��&d(���x��V \��Ln9��RK�s�ZB�7C�7��(!��^O��z��#���mʳ6�:	���+�ی5=DW�4-����g��㋞��	�ݞD Q�B3Ę�R��Ҿ��F%��v�/n��i���2$0[:k�ކ^2�t�)"�Qm��|���Q��9�%���~9$�3�/���W	�_%�o�<�,0εr̃\~����d7��Ez"�_� �=x_�e����	���H���7�!N���Ζ|�0��9��]��	��$>T��w�K@�?�{���~�:��錄��fa�F8G��d�g�-�|�MLMH>|��<���
��� �0�8��S��#�����xK �&Y.�%%��j����୒�[�'
��<�߳�p��~(��$v���
��\�+��|y��+���
;�?�:z)[�:N>�,�TIM����=d�怅��d|�Ư��!b�102�	� *9�#n3���/�G���hy��2d��/F~�5ەm;����R ����Y���s�a|�8���/y���'|V�>������W ǟ�_�-�d�����O���&V��u��Tof��D�kRR��(��H0k9K�U���]�p%69?�w�]����t��a:W������[�WK�Q�s#�{���N'��|p�a�RȃY����=D�5UDa^�nj����Eb��R�3��	����.���f�.`S�t�rjgq=��ifO"��q��s�i"������Sxչ�ι#9`��m*�V.�����de��Z����l�%q�H(xؒI�v�9Sʾ)B�I���۽���Xn��V���X��=��l6>��ˏ|{̗ꨘ��˩�	-oq�%ݯCM�>|&)T��x+�<�,�x�鈋k�P���t��ěAF��8l�2/�P>��j�;%vBU�Ϸ;�H��'����S���z-A��N�)�װ�|���'�#;r������Ӽ?��H�o���;ٵɳ�6M�mغ}kSrlv2��<*w܈�cv	�)eM�Z?���>LwWG�|9��-��pe�MWY�����Q�Sn ���9���'�s�h��P����T��[�n�5�
�1����}D�Q�IA�#����h�y�8k�^��.�(��o�� s>Z���t-�)��Lc��E���?��2�x�\H��4�/�*��_��dX���4����DĢ�M}�1!�*1g��s�n�Jh(��D��j�|M�d3B���dc.�{�����I�)%�������6m��u�
?�LPrt�!���3_D���
~��l����5-a��y#�>��6:'���p����N.W��Mo���I��ɢ�w?3��\65ǃ��}\4:�8kFL���J��������V<��af �QNb1?�nT)�$�
��o�����
����8DVX�D�{4��5��MD8����ׅ`z�B���#���&���Cs��B���ۆ�C����հ����F��UQ����W����жez�靫7U�Zۦ���n�s%���Sږ��i����#�1�g�ű���sL��+`qӲF���8�kz���?v�$�Rљ�S �_T���%�С|T�����"$��{ݒ��7N��g=*���L�;*v�!#�ߦ�`g~���F3��-,��L]��<�)Ud��{4�G�VK��^�=� �Z��*@�HM�7�@��S��ʮ������:��xK�8�$M-���S�C8uϩ�%�&�/8m��3�YB�*�? ;$�b�Q��2z�!��"����^�3�q�+<��@!"ݨ(���:�7�����%@݀�k�7�} m�����T��B�@v�D��ȅ���΋̔RC�lw�����7�ʗdA�wbQqr@�L��+Wy�"M+��j����\h�
4�AiI(����e�ݟp��������6tJd�t�B㺍}�R��w�<&���&���ՙ|O�'�����c�ƽ���e�n�¿�o麒]���F�&���z������WY
�t���.�5�a��6��@�5��Q<�9��	P���Z��"̾ר0���Kֻ�/tt����'4N?etM\:�{ϰ��ԅ_�7�6�lx�sK9��PD!���
 R�����YXB�A�$w��Oٸ�8_���p[d^բC���P�o�4ր�t�v~�/k ����u��E;2�����G`�4��<)@P�\����:k���(z<� I<z�r���� �a )�9�����NE���n	V.���Xj�je�PN7_��z_�+��9�s�����	|'3����+��v1J�b|¦��K��j_�,\ $���#L������ɦ����Ѽ�ݏ�U}R�!ǟ�1�o�=�MI_-�*������w=i���D7��$aף���e�����Yi�<r|,��D|z�Y���i��X����K�8$�N:�Q�-����u����O�<����"�(���7u����s&J�m�b�3ˀ�ܖLE=]�ߠ���J�b�?]P~8k�&� �cӞ��⠛m4���ztJ^��u�q�h�n�Q��p�c�ҙU���]o������� �~���ũ�qj�� l��^r�摑� �����e����`��j��~q�?1���0�����k��W��	�/���W�J왰�^&+�2s��ޮ����[��a���=�u�������^�"W�;�P�z�udj|wF����0e��.;��x�$�0.m�H_.r����	vp��d�*�.j��*�Nb���;�խRU~��'�0���d�C+��"�P;o�E��B\�l_���N
m���ܿM���M��O��3�'�W�rȖ��ز�������btP%���#��t6����!y��_��4��x�L{���� �ow�U��-���[�����-�q=v��hmX��^��Ǚ�'D~Zt%��X�9tyiY:��3��� �� ��2�Bϸ8�kV{�TnJ� �fv�c���b�-�{��֣�_��\1�9�_Jh��j�P"��X�e��n�le�ZX�_���:n�K�z����X�.u6�N��U='�<TOa}�@Z������W.E�d�I��+�y��g&�x̰7�Ν�i�����`��柧�M�ꆘ���t�q��Z+�a4�l��f�q��~v��;9���$���)ݦ"JZ��1�wZO.���_ST�,i��z"��M��t|<��-��2��g��9��^�<@U��$�T� a������6P�Ɨ}T�s���6@�����"@�����xnoc�-��Q ��Y���g>8kFf!-ت����!���TE�*A�Ґ�k�k�ۼT,ĥ#<p��D'�+�U�jm$�r���R�!�o<�9����0�8�Ѽ�� �K��B�J�&Gm>Ft�[�9u{
"�����!I?������թ���Ci~2�,t�sr	�#�4F5�o����$^�s<p-@�Zj�4���z���s�kEk�,��YЖ���>V�Bt�%�z�%yh��jp��f'=AhC�M�	����Y�ը�W��m/Ѩy�Wy�5�%�U��|~���V���⃷���u��C�|Dt��ݤn�
u[�l �����w.��� !f���@�s��tsD�5v�-3�~��zG��D-/u�Mh{��dZe��`�N�F��/�x�n+ G�Iۏ������%ȁu�N���Q��h��sv$�̽��p$��?-�࠙4�d�}$+�q�]���n�/����.�/w���8ڐ�'�s"QSTn���5}_�k���D�����~Nޥ�j|�硛�=�~�HA�;��GP'�	�}<�.�1�E%1�E���B���LA��UIb:��ld���)i" �R�.@�;=�ES���ř����]s����\����z�׀�[!#Vi���a+W����Z
=�Nf�fl�l	�o�l�WMG��<C�J9`���8נ4�ez0H��=dB�p�C'u�k�JX_4�E��l�s���ae�p���n��kD	���&�s�ݝ��ǅ�Bƚ��{'�����S��1���
���4����Z8���&��7G֎���M�N�Zn�vh�a74�z�w�QR^ӣ�`b=�N�ZH\"��ԅ��c�ʑ�ne��G.t�sȯ��c�9r �bOJ�:5�vg��?��;(}谐6���(TΊ��t*��l�8�B�Џ��1�1�p���o�7r:�r=衅(��4�Gu��`��:�����t8��3�"�g�f���4�(-)���եYD�ULL�+��N^Kб��<��;o��)K���@�t���ʞ��!~"��/@�?�T���@0,ɉ�?�����LPOP���HCGkZ��ڞ�gQ� ��b��8	�(�2P<�n;d�c�
8���9�-����T��.�~��0M�-�����G�k����Œ�q���.�ƹR�;�(�`�fc'��kuJ8�:]��٥l�iW��H�FD���g}�[��u�8p�@W���G%Ad�������Q0<q�8Qb\zNlz����ƪ#5�B2hJ�fݙ�
��*yqe0���;��j����VR%���'}�͡�� ���Ks뱛��%Ln>���e�М;���׺'k-p�x�1���W�",j��{�������˭��u�NT4V��S��A)�Dُ#�z2 �-=�ta�<*~I[#��	'������ܬ����\Y�hJ�(��<�E�-���$�܂��a`"�c��K�/�~k�Y�Ҍ]�~�NO/�Z��5&����$�Mn�z*����I��#QپY"W�k��ӵ�e�H
0����X)@S_f[<ő��D=�Λ�q�xW ?�|>P2(-�]SȖ+���^�JR D���K�����H�~�=�Yw�/��S�_���Xz����yx��8y>�����<��f�u�K+����'�I��&��pg(�lwIE�&��'C�����3�ތ�j��lB�!�� 8�CQ)�F���?fBu��-!�Ϊ��&g��k0���fjWz�F��%�\#h��`�9=�]�\�a�:%�-Ak�5T<����N.���)�����C����k���y�d�#7�H������L=����|��o�p��M�LRt����%��|c-[R�`�Ф$��dY�CEeH��p���h�h�Buκ�g� ��P5Z{珺�=��&�<�䟛�t��6(e�y�f��^��;!�)O�Q@�{�s�zW�0�-s�(A���(�%1]g���z��~��'r5��xX��&a1�^i����d87��ճ#�Ȍ�P\[�飯�c'�2���5en��T6�v��!�^Yy������=�2�@�����U���
D�Xԏ|��;�:������U���{�>+�y?�W\�>�1��� ���E���4��IK��5�l3�h����Z�/
	���hjm����L�A��m�l�g7��ly�x�L=,��*����� 5�ؓ�b0p:��`an� �+=�|��W ����j�n�r��g��Nrd�Yd�iy��M��4y�E��v��#x�&�/܌�ګ	�!w�>��<�N_}�g7s������X�Z�i]�|8������sQ�KG���\AG�m<��a�K"+A�"�C��Vx���
ߕ`�'���s|&��>F-
��A�
{�Oۑ��n[��m�é�W�#^�XA��f�T��
g	p�cwh�~�_@����J�&&^�1/I6Ȇ��Ȇ��MA�P��} s����(�tG���C���<b��`$�Ԉe�?���h���D����d�=�%��R���ϔ/p,�� $����y��)h��@g��Ʈ��ڪ��G��g����G��dIF+;�y��y9ܒ���>l�	o#���r���=h1DF����U�F2K`�ܻ"Z�ʻ\e~i8y�K2��&�����}���꨾ʒqUQX%�@�6"�$#��j���B�H�8�v�3r2�p���~�,|m��E*^�UK��P���/&����D9����ޜ�	EE�k��C���tb�����<��2Z��:�����4��Jվ��lI�81����l^�d>q��gR@��8��]HpI�
�_I^M5Ad�#�m�q�(�y����Z��Vp;WiC�1���g2l;�R�>e��tqʹ�yn1��jV�v�������'���_��a����Ŏr/���
�=������_���UB	�I	��e���K���'?�6�-��d�M�2��G�nL��P��仺�&�e**yҥ�B�`n�]v%R��x�Z{�~u�c1�	��������b�l�nG3��o�u������*����i�4�4Բ�RD�xW�<\�	,n��vm��@_HU'���$�����`�Aq�c��)�a���d@+s�= ��CqY��9�s$L��2�UǞ��o��a�(Ej\CN��������H�J�o���9&y��ٲ���+$B�E~#"A��Dn��|�V��
���<�2��݂�+v>�N#d�Ч�Rh�w�% �M�k��lͲV�E,�U��B�����|ti�r>�.�Xxw���7$�>.�ۼ��/[�)�Q_"��@�����o/"�8D��*zI�CgT�K�� �h�g�%�8/6#+6��ZAU:GH=!�L� 'ä_x_643�{������V��~�m���g_����6B)��׏���,�̏�M�7.G�N�\z��w2�G�]��c=	�K���h߂����Sm��Ea"�B�u��#�g�0�<G�aD���㛏W�oM�z������X���&�>���i�k�n�HT�����*��S�z��ߖ��_���14�t����Uw9�Z�_k^}R�#N4٥@����$��8j��� ���^X*O���z�_w_��p:4C/b�,Y�V������"3/��K�/{(�O6NF��{���̃��C~8�s\�*0l�DN�u�_�aLi+�����\���z�
Gm����mIh�����X�`Q��z�d�r��u����*@u�xA��;��~��Q�G����QVsJnCX�����&����I�&�������q�{\IǄH̑6Hғ"��N�aOO�8<Za���{|{�+n��|�z,fTq'�S�a9��Ղ�u�+tD\n�N�N�+���USgđ�$�M]>+���@������H�X����qFr|�K}:�a��}�@2��Q`�����K{�}�
�'���@�ߖ��6
(��޷,��5x}p�JpVg�� fp/۵$�ȸ�~��:�˸��������(<�a��OPH7��Қ�q��v�+G��E�=� u�'{��ڼ�1k������5XN�y�� e��X;���_�Z��qu�0�rP�!�T6K�D|���D�T]�S�:K�fĄh��r�;<�L�/}~ky��$8�����C 2��j�s�%�xA7��#�V \���Dd#����%=%�@�n�nߕ�J2�Y�4�h|$�c�۳�u���q��<�^�sX
�lO�2(6�>����w�wZ��߇P��$h��S�/Wf��<�����s�M��#�4[�ebNΉ4��˶��`,v��S�䅬�#��������v ��$�B�^��M2�\��3�4[�]o�����5n�y�Dw�g����������;�C\�.|��R �� ���A��S}B�LO���OoY���f�q͛��vy��wU�d�	�i52�G��,���q
v��o�p��������Ļ���k�u� l�}Rfښ�T~���?0�sO׭�7�\�Sna(#V�x���R����D�@��r�V
��[��$?�,o��}�A�	T�k��奵9g�g5���%��o�B==D͙J�?yc{a66#D���-�4��2�&l���5���=�s(�9��Ð��C�,j?��j�3��L���42�G�����|���P�Z�O����j���1p������=�rv��̏@e�/���o�G���e:���
R�҅��Ԅ�>Z��Q� w!ێ���6"h������Dg�V��&�Dx�E=�M�<>�g�&��=.-�1��i_��+�|�r=C5l͔o���r�������1�L�Z�������+&;KsB>C\�n�P��Fr]?�������@��Ol��5�Ќ�����2>h��(|-����d���)c��ԛ�2�a����rH�I��C@QUi��yf"z)v&,<$?˴hy�}O�)Gep�x{"<j}�S���rB	9Y{������6�+�r#�@��_��N��`N����x���܇�Pu"�G��;Fe Y�>5���"}��� �6���i|����FX5{�ѭ8K��,�D-����r���iW��I���'e��+Ż�Ark�-�{_Q�	!�2���3������йX��6�ZI��RvM�En0��/F�Rd{��8�4�4����2¦��BT�#��D_��M�䲕����tB��C�"0=�߿0�/��� j}��̷��탈�,��`/��b"4Es"�?��F�Ĭc��R=�A
�q�n-f*P��	��bR��7�X�&.ֹr>*��[��%I��e!��?%�@�+%�t@���HH7��P�C��[���������K	�77�e�	�_]�X<��d��o��>��~��qm?�n[u����h5�4	���8�P�td����VhX��po�&y7�!�1�l�J�ѵ~C���}8<"AR����B�fU�e�~ ���h�R��(�/�
>E�nz|�4�F۞��$�pp+��	q�TTqFW6#�O.	�A$���qF������)�L���ı����r�J�ř����K=|��.���X|ל������/8%���Z��;}j@a3�)��²>5�Nv���91�c��&�V��n*����ݷU(���MQᒅ#fR�����Z��� �����L˞��!=�yM<3�V%v4�ը��%^�& }��7?��U]���q�|)h�M���zrBMa9�Q��rh�������t�fi6���l܁�1q�rk�Te����<����_:@�Kn�Z��9�:QK��Z��������)}ߑf�1X�f�����h��}y�b��N�`����2)�g-Ѵ�@��toI�K��{((�R-W������a�F�v�[��`�[�֮9����v��F�[�"ը��v��Ҩ$I�*y�H�m�|�]����F�Z���j���j�2L���]>�Iѯ^S$�?�9�*�\a�<z�)�Km���v�$CI&�#�4;貳�ڝ��Ο����2R�v"�c�fq߯ZG����[�c����}�Zr�9�]sTς
���������L�PÃ��;^��
Zcal���_��n���1�p?��kϡa´G�[��`�Ί�)'����L�;kǙP���C݅P�H�t��R����H���7!�|PY&�9���҄E�u�B�24g� ��Ii����� v�B�.����O����q
m�$	$�jS/+g�:<;;���$�7+v�p��?+Fdάg�BWdv�]f��}J�n�̌��ҷ�L�2+����-�{����Ih̶
�5br~�K���H��HΡ�6���箙�oLt=�@nƝ��G�+0���@��5����ū�	#�D⑀b�#��Ve���^��zSa`҉��q�PA��cƥ��m��8�`�m�d�]�>�]�1�3�c̑|atִ	)����Nb�K��z��]PO��f���m�i���4/�q̼c��X���
D��d��|��nZ_!�>x�§L4E�r/�rf�L��u��Ϊ�۽��x�s��,�-�2��=T������i��_�#{�B,Ú��l�`�����^�UR�fin��va�_l��yMl�����2=W���Qḃ�/�p�-%3`r�Puz'���B.�_m�_X���hK^���T�R���A)�C�&$4K��5cC]��+!df��r�w�'2��q�hQ���j���a1(����g�-��('�9�D؂F��m3�^:��]�=�6��]�^P����#&k�%�<9.��?-���@Y�3�g�>��E؅�����1z��kTQ�l�^;�Ӿ���4��;�e�$�?G]HkLF��񒮍u�(xn����Ǐ�L>9����G��w�$X��/��Vbd䕀�[ `'�� T�jg���Ĉs�a�qٿ�lpK�[2��,-۹C��'Q1�����
���8�:��# ��J�a穓�.��ʒ��Qo0ɵ">Ѥe9� �M3�	%�S��Du[/6@0�[��L.����*��7k��j��_�@Z�O9�j^���ǰ�Sf��XZ_���k�Җ{�&��u9�������1�?R��?��t8,Sb�h*>� �G��rP�w�)ϴ�y�we�Ft����f��}��bI�ά��{�VM
�g�țE� ��{��b(-������1Q�U��*�x�4 UXS��lx��NѬ�"�;��	�[e�DM	<���1I�vI�#�U���䍀e�\K�,��z>�
r9�e͇K�?,ġb�Y���/�c��rT`��ǺJ��s�	+�?T��>�>��/��@|3�a�{Ó�8|�q��:`
���_�F�3��&"���PZ>
Zd�!�4J�04����.��M���E=��aq�تg������1���q�1��7�U�0���/�D��z� ��+EΑ
 �~7.3�]J�FxWՁ���/>�!te��+B���Mc���)���_A�NdQ�l�y���	GDJ���T�1�J�(������"�U(;#V�)���W/0t��6�(�Y,�}b�I�eݻ���4�����d�Re�>���C����t�~�98�#TM'|eo@��Z��i	(��{ǥ��}`u߀D�������`��xZ�ձ����j0L��"��κ��!���ocV��+�O4���Ȅ���Dh��B�_{�F=�T*)�s]O���|3am|f<��7A��w2H��(�gY4�fJ���q?~h�W���{�o<�lt�F�P�O`�`\��R���+TwVN�dl�!ov1��<����y�'l��c[BT
�i�Ҥ}�3�lg�f(�[��3�g;E��yH ��h�:R���gN�CX>i(3It�z @����i�h?� �Ѯ���]��=��Q6������}�K�M�ώΙ�Ց�����L#חe1'�� ���O%'6�G��3�@�N�����C\��er����?�֪��p��<�Ssן��Cl�ր��G�����05t������SKH%_|FY4셄Dt�qTO�p�~�7`^}��6qx�hA�NO�c��@���)j�G���������X���{;6��a���V�����;45��b�$_X����6����o�l7�pp�X�V?UTA��푼NR=�-�G<�կ��]�3[�em�?E	��f�Zn�����˯�T/��i��W2u��r4h&�?�O�?��*���3�i�N4�x��TW#���l�k���[bLL{��z{�E��Qv�d�'K3�`[f�6�>PX�m��뜃��a��b������I,_��`�J��z>��R��)���C���?�#\g%k����D��=�d:I0|,�䑽Dy�Κ_7A�6�yݭ(lA�����9l<���O$�l��q);ej&�,s���MB��u4M.4?�Y���0����A˖�q�:���?�IN�ش"���ד�1�Fb��W�j����םV�TZ��;H�o��hߙ�W��0�9c)�D�*s�Xl����y�.л�as	�7yH�lQ�<_uE��i��o���J��aX���f�\��˩:T�\�a`M�g�mG}5g��}1)=��yL�4n냬��k�-~�.Hi��0��V�q�,���e��DViަ:��H�};eh��HQ���"2�Eͬ��o<�L\�gr��%"D�aZ��ki���8�9��U����f�H�R��KvτZjVP#�X�݉4�J�J]�~4�� l!�<�?��z�����<x��t"���O<?3;��V��\+�j�=�Ge&N6}i�V	{�,���N�(�LMfA�b��������5���#��.��;J�ab�*��Ã�＂���c�L<tDQ��	N�IU%���d�!����<�eӘ3���AZPz �u�
����2���&8	���t����� "q�e���KՋyZl%+�ww(ٶj�R�²H�����M���3��՞A�e��r蜍[0�S�O�o�k�:�%{<$����r�|�/�x�1����s"�����L��^g�����T��A�3Y;��O��s�@2������{ל��[�/I�&&�th���28G��m �pSm=�nR��CT�" �?�P�~��"�Ǣ�Oxkrz��?�g"'�!Y�nv�Y=]z��)<���b��X�O�s�#����f��j�L�w�iA�{Jލ�������-2-�?\h�E1m({�_��pĩ?��.a����OJ���$�Z��*`'k�/r��1p)�{Y/��H�+��@ޝ�����3$��MY�yc2(@o�~Q˚S�3�o�vr�v�%D�I��:[3qԑV�I-b��d�*��:������� ]~��ΰ%_���oܥ+����m"p���8�'����B��78p��6��X�ٔB����љ��KG��s�?�&˕"1,0ͫ�+q@��Gb 'kZͬ�D���J��s�W�,;]\�q�F����O({&	ͅ�A���h<��'�~8�.�Y��D��9����񡬾�����3~�C7�E�D��he6m��:�%3-����qix�M֝:1�#�1ԥ[|�V�J���D��Bt6d8F��!�h��lN� �
j8�W��d���O��L�**�sx#�gB����l�m��^��Qo�f�I���i*F�*��۬ ~r��6�y����$��;\B�r�_;�mC[����6y��f�F����6��a�4����h߷��װ,����-������+RՉ�L�o`R���ޖ��\3���������>1`��Z�U��>P�������;xb���!�=�e�!������j֮tYJʻ��H�0o	9���k|G)v0�A�� l�W4�KBF�f�gS�u�9��]�h� D����A�����\��6N}�b2+����߂Sײsq��j~#Ie�'��BTh��U�2�Qz���X��5��G}w�,��6^�_@��!�/�h��P������u� �ҳ�|�$���NyI���t�@�,Z���?�D���pw�0���05���]�*���W&,tФ�2�`Ք�
_<�U�¨�ҵ�z�,H��Ѹ?�(�X;� �n�Qù������Q�Ě�tn��Si�~�B��8��(��+��hh��E�'�ױ�D*�ڶhpD �� �+Dj1�������]iZ7��<�H���F��&���Ly�b)�G1h��`|�T�ey��?�< �
�v�V��A�' ���{
��*޹�J��y|�_h[���L�K�nNE��^���c�����+������B7Iu4��1hڪ�A��nߏט<�0_F'z����̮M~Z����w"uM\�Ӽ�&���e{��S�sl-��Y隼�t���T��
wm�C�����I����9y�A��<���GWA�s���OSj<���a�'�'�)������}�ի�� �x�SO���د-�
�pSد��b�:t,�Hi��Z���1`!���j!�q���]��*�Z��'�o�(G4�u�N���:׺�&Y��6u�:�,�����6�k[g,<'~
�
��T�wmF���3��`o�D�"��t������V�"���ɣZ����1�w�����r_�o�>�]"Y���	d��d'O��6�0�mV0)�qp�o5�;ǡ�^y����9�������O�Pn%M���3�^L��g9_�Pkg���$�d�Ѫ)/��{����gB��O(�V������B�'	%���ڴ*Yo`���=o(�9f9��ց�.<��,k��fȰ�`ǥ�j�L�b�����h������8v��*$G��[ȴ�[�w�Ai��u�lnc�吇2�ɸ�g�Z�<W���5e�Zq�S��I�z�������Z�b	���%r��!�8�㼃v͟w�eU`���#ҍv�u�%��GVg���W.e˟�n{Zz�6���&���lM��Qy@�fr����'2դh�3cv
w> s���9Y�P�&}����~�o, ;HL��]�۶`P{|�Sfs���q���>�;\l�dļUnH��ӟ�wE���jx�#���9�����2�I�/$����:�
�>>��= ��5�(�O���):�c-��m|���*e����Ek�iɨ
��U�2���~�d$l�d%�pp$���߯�UOsX�-&G�:_y������;�09��q=ع�Z��8�\�7R��nȋ�����;���fC�����u,��KL�)�yXX�FU)5���S't��G���8cO�� ��������W�`�_�V�z�r\�9�ad�̜�n�do�q�w*��	��^ռ���4=�c�a�'�>����PvW�س�}�+����5�9
����N������������J�~ecd!��e������j�j �`�\C/*�BSux�z4�8[l.�'��W���n11�S8ޅt.�p1��W���;���
����EV��a��b�%n��NP(�����Y��?��	�qLTQm�q�)�4�
����Z
�cv�¨i��r�m�8��P��s��CZ=H:���+Oi��CZ�����.�SO��
�l�^���ðQ�z �����w��D����k�pೇ/��`��O����X���v���ۦ������O���`L�Qɥ��c� ��&K�@8�U�]��J�;�Zƛ�v��#�]��
F����j|7W$H&8ٗQ1&Ά��.�p��7 t%rF!1t�W���d��ܼ����O3��SH�UF���U��k���������ֿ>n�qUC��-/i/.˹�c���WY��5��^�A`�?���a��[m7a���UA8ǈ�Y��t�����iǗ%%>�2Ii\�w�Z ����\��Ҹ~�9���_,������@�n8㨪�����������S�Bac��ʊ���sBN��b:$ ������J����C��9��R4�!.&]����r%Oͽp���m�ġ}o_�-Ku�t�O�zP�ז3�CԔ���x���u��"����]�n`�1�i�Ot�ۗg�4ò����u	���!)œ��d�q�����/��0l�����Xu#���2&5X���b��+~�λnd�	X��!�C��P��5�o��x�`�b��Ta�l�:w�;AԩS��+r�F��Q�����:+�۳�^�
YurB�͡x �(�7�%�(��a���JX�#���e�F'I�st�A}�ꃱ-��#5ޫf�V!�k~%��B�ט���
r�K�wc3%җ�W�X=_����at@�#�
?J;p��~y�z����!����*?��@���wDE^��ϗ���& �QY�O�e?�1�q�N�y��>�u�b��Q#zb�Gڃ�^��z!kvx��ܶ�L%,Д�a��Ff�r�ͷ/�3\r(6hS?cNq:#o��)$;�=ˮB�~)�h.� Y�6`٫�8��������_P�*3'Dd
%H��:[]�S~���\�e���uӔd����9�
J�A�;�6K�bh&4�"(�:�-ָ���4z���g)R��ߠDI��J��:����X�0�q���b�������F:Y�2�`C3O�+������I����P�����w�9�g�R��p����m�1��܃��L� �{�D-��b��KE�L�<(�X���Щ8��
V�ۦ�xk��z�Yr�w��RD��C |:W`�>ůڮ�O�Bj�К�G�Y��X�:Wt�nBa���p�,����忍qyT����A�|}�z�Ů<���@�����K�g�`t5��1:�1ݳ�fQ���>������dF��ݿ���Sh����Գ�y0[�a�z�^�o�SW\��AVo� $)x������n�t�6ĕ:XE���@a:���t�B����]�d��5�u��i�N����$2�$����U��SU�;�?E;�ͺ3qtT���Ӛ�W>:�Ђ+Ms��5�G�$͕�M�a����g$9�*l����#�t�.v�-�~$>ȈT���g�lu�\I;��(OXcH�@���T��x��]�J(�AJ�G_��!��������4í��"MV���������%F��B����c!���:�q�,��C�g�� G�A���u�� 6��G{�_�_�*w�k�\�r!X�+5�]L�_�&]�8�'S��Ӣ˝�w
�{g��80��J���a$)��&��䉰׊��7�a ���Y�I����!}� �騬[���j�K?���2I(G�25\G`��b������pNf�"��~We&�y�ң��5h�D����M�~{н��w�d���{��!������͟J��fħ��K�g�splq0�����/���Gm`:m��b��`č�^iOn���I�ϭgu����H
c��}y 9�����_gF�k#�)^Ъ���:����\�G{����ZC�uJĂq�	������9��j�_���+����� X�� �w�3�YS5�#�`�r�=��$�N	�L��#��t.�+�0)^���Gg���hP�fzhgĬ��%r�:����X��&��'!�T��4Ou����������y2އ`��y�N�9GG6K5� �AB,�Q� �ч���A`������?�J��xs3�7n�b�X;�Ȃ�n�n�{x�!.+#��
�(HϜ��
b�6:��X�?���a-UP�c�Gl�Ǡ{o�If���>��%7�����Y�FV�KX���O�)��o��  B�k����=��%���	ÿ��������#��)�K�?_�Ω��4����/�[U����1"+��lRU
�_7=@��a�̶驰�� ���R,����"7�z
+jQ�U���6t�ݍ����
C��	� �Օ��M@w�B4��i?~w�yG�r ��=	�[����֟�z�'�r�K�}����Z�^L�.4FIw��,�M�0��%������+����EX�XWe,7��we��
Xvޫ����c�wҭ����z�Ć��I��f����=m~�ˑ�6LK���
8c�!���'�W���"(I&Z�-<�ط�&��AH�T1,�D�����vH�_�ޑ ����Τ��/��f����ѝ�������"N���$J'�!ٮ�a*v: �+��π�����r��������v��LQ���a���'>��V�?�� R%7�!�>$Y?ا}�L�J����g�h�1�\9ʗ�Nx��z��{x�r�(��,�yz��]����ŗ�ʥ^�=-�������ǿ��q�{�*�i��g�w�ZH �f]�Dw-s��H y_^�bUB��j���!fr�kq�c�j�]X�1f'��o�ܜ������@2g�r�bs#�0&�vS��QҔ�+(4��9�`��&ŤN`R�F��'��7H0^²k�d`=���t�9 ��8�9.�Lك�K���ruY����e�3�"�Lܳ�ް���ɔV�\DXl������2fV:b��L�)%�R���{��T�[���=��~���w��t ��H��mI�:���1Q������M���ȦS �B�T�.^���Ɇ��Y2Of�X��-�zA�D2�-<eF&�Q�j���V�w�꾂��[�DR���O�P��u���3QZ���]�A
��
sL	�"� ~�(��Zf������_�Qa�Gi�?����C�S!M�9�aS@b��_�7g�xw|*gx���
w�v�2ͭ�Ǔm�d�ka�"Pݙ9e3��!��rw�k���WE�Ȍ*�,>����w�]G�){D���Q�t���� ��a�G�YZ�?Qr
��� ��N�́,� k� ��v�DFTz�B��8�J�U1���6aCݿ�!ˏ$��nj��x�ǝPJ�n�Ϯ��t�O+D��#Pٿ���h&�T^)�h3cu��Q��C�'��<Da*5T�i�cY?�*�L���d�s&,"5��s!['�����l1VJ0�������O�j��V!WF�12�:y���UNH(p��NL�����*��L�g��R]��xN�8����%S�#*�N�A��6b�0b�dDFA�Н����6I���(�'N@@�h��D�β�jp����ȑ��u5c{ ��L�ڗ�H��9b�xm�K 8�����&^����I���/]�Z@ql���g,6��>�&'⯁D�L���N{��D��x{x�Tc��zr�T1�c�=��|�8��_`&�,����e�j�>�9r���V_%�K np��`�Y��������� ��@1At��^�z���Uw��;䖊�ћ�!߯��N�U�<��֗���ϫ%�ssj6[H��a��/���OH#�E/�W��*��C�垮��P�?@�m�:<��ez�m�eZ�(����}`d�z���jֵ��%nZ�e�QFHG%-��I��������U���=��/����e��c�FO@2瓌s �7�_��۳�F0�}@�/��Z 3���ǗGoܺ҂7XCOkL$�P&�p��'Zx��*�J'�rn���S���{3j4�i|����1_��4�e19[&H�<��vG���3L��e�.Q��v�����4Dݶ�|$K�V��_�wfkQ}n��+oX�|!�M�|��ǝ*��YAL�>�˞E��U{Ti��:0Pn�:�%�tƒ�0��R���_v
xC=�$�k���j��!�o�
��b���W>�Һp8E��@�v�����������m�>�2Ђ����N�H،k�����D�W�W���i�N �a�dj�������]y�d���"���)�[���QҔg���	��S�yS~ND�s�۝ꏒ�2L7s�ts��G��(�Q�#;�sN���;�⢽����
~J���c��Sd��2~b��#�]/����1�wJ�G��j�����X�I�E�kb���`"�}{+���9�e��'�oN��~�"{���NZ����L���,q1��a��o$F ���(��]@�˨�s��:A�Ŝ3�4mWXL�M:1b�`�I	�����48�Ƀ�(���-C�O�����
;���c4�!x�%��[�R�Pڽ�ik���y�_F�~0�	�0A�zդ�[Vh59ּ}˝f���ǐ�����U�����ikh�	�>���
�ϻ�T����1�J8d��N՞80�:�=��?�;CtT)��F��"�:X�A!7���M>'y�0�E�	�R��w���:��B<�����	3������p��&uW���1�h� ��%��f�D���>\Ѽ��?��O5{WK瞕�.XtO�����1��_�V�A&��'��.�xA��.fs���\s$;r&י̝|�:Rd4���a�dT~��)��l�z����sXV�;� aץ�U�UJ���}"P!�{�z�A�A�,Z��`>��P�=�m ��~q�[jr3��F���3�ߘG��R��[�O��c$0�Ze�ƴr<(\_-q�E�^q
�CE�����B.�]�P����fI�u)�p��\�'��S�hzsX���]b��9�\E5�n��]��U���nX�)L�dY��r�<�AD�M��;�C!� Jbmd]$����$�s)m ?�B�\:�A�㗁k�v�ґ�(�DM��x?�������,�h'㦴�'~���a�H�5~����rP	�8jg�AP9�f ��>U�8�T%�XjpN���0i��=AN�xfjP��7@A�Ʋ�~��2�wgu�Ҫܰ̀/�
_u�|EQ�?�<���8�6|��X��7���Ѣ�4�5W�6k�)E2'xyO��77�,����(�_̓7��U[[�$-.
5Epk4��w��ԄQ������P�gt�M�3�
bGR%Lf��z֥�Fշ�L
�u`��v_6[�e7`A�?���~)���[X\+�����K�ϼ$�
���	�$��������P���hl���aqhb�f䜔��~}B���+%h}ǿS��nö��w�@L��:O0�
?q�[-��e�~���M��2\�n��):�ExAj�i!�c$>G��k���"Y+zC��k�gl�&�?S�!�Ə�{��*�f�%��hE|��c�(�KS2�՘�i�"����m^ݡ|`p��=�%�e~$ƪ���e�!��-8L�AK��/o��3Z�'�JJ�A�Q�$�����hg��{�� 7�0����ﴼ�"����@�Ȳ�~V��MܩP���:��'7�!fW�`1av8��+0��?ά�>b�Ug�m ���%�� 8-5dϔ����A��n2 v�Y4�}zh, ��L67m_�|3I�rLnȠ���w�}���N�-��l�HXn�b��s����0��j 6c�q�}�{��A���lT��ɸԛ�u~�ҍ����hR����YTs<%\jȦ�8q�T���P��[�٧��x�ʒ��4��rD�?���{5���6~r�h'��ԇ��[P���sH��,�G�pX��R����'�98�}͗\�&��I�f^S-�����܀M�`�fN:X��Sd^c���\��ůBd(*�l�N�df���]��by������Z�Z��+�۷s'F�֐�y����y&o�syn-�Xu^4)�r-/��2�p<w��� ���-���ny:U���ˮ���:�w禬o,A8�	4jT.s��d�}a��ڇ ����п� ��8����F��ߝ?�`�@gR�G$�!��QQI|p�R)�C��'Q�E/�ـEH���r	l�u�D3�3Cʾ� ��J�Q����B	�;4��7�I��	b�:��R?a~�	wܡ}[Eλ��Ȼ��!���h�ٻy���L�AJ $MBM|�]��Lg��  ���R	U�/|�������k袋\�lp��	�fW��
Ȅ�qh񖴞F���Wsi� �9&��e�~a#��l�!wS�"^D��"8�N�x��c����זֵ�^m�j�"feE��d\&��(qK��Yt�L:Wi_׾�\����ȋ�[�0lؿ��*�����^w0���b��+*)aU�p�@Pڐ_�����J��G�*0�L��-Ҙ7�T�Hk�,!]1�|�z��'5���,�X~���`��N;M�\m�P�����8��<��a?�a.�x��\��n�
N��u�et�&i��0$���ޱ���@j��yP�hEzπ�okh6+`���}8�o�q���P͆�2�t�9�͓hQN�S�aC,}a���,�pq
�����+� Y��|��g��#�@��/�����-�HB���T�
h7~o��I�#n�+Wi�:�2��H�&@�j�zM­
b-���h���=%�ǶG����ctp��	b��~�T��-u�G���X��;ǀZ&����6!;N�,N�`�L�;��:����mҁ= �p��2X���J����؄x����r��J�l��'�>M���B)�m�u�!~��%��T#i}���u:���-M��`�B4v��Ͼe�!Pv�<n/��x
zҭ���4�~D�bVU��N\%����DV�~r��.ǽ!�c��\�Eն�?	J��^��;p�����|8���C�L0�@��D�k�B�B�����6:u�rŵ��Q峁}4����Z`��f�ST5�d��D�m�%�[���S2���Ăߍ�	g��'F��|��@�/xM�� ���+8�b�?G�.����Z���!ы��S�D��;Ԯ��2�da52��ٍ�]Շ�I�\�>U0��vR�������3T�Y>��w��¬�5��ŷ����%�L硜Gey�	��������^�;��B�W�z�[��U� �GՀ�&�k����֏��L�dX�s�3�ő����ΖeI�0F
���8g��	��aܼ�������=!ړb|��2
\����b����@�`����9�g��s�6Ѕ�"JY_�)	����H	q63�"f���r	Ɂ�� ��5.6N�<�l*�Tp�&w�� �b0u�b4t�Nן6��$w����,|�d��:����(X���1�\Xl%�r�ߕ���Eh�Y�s�����(l�mPRې�(�:��ȸ�'!��kۥ�& ����L�6�O��zS�����#5���Ù�V\��[M!_u� ]v�XuM8�p�]*��V���L0x�W�Q^����f��c���Dp,�!��|�����N���4�$�*�=K@�>R�~D`��-E�U��zC��Q�q%�ժy>��XYV��Xa���[Gb �f��zZ�;��8YKzז�����ԃx�ǟ�<�*v75��:�d����Pe�'��}�rL���?��b$.`}�9PD�#z�\Ӆ����"��zH5��gy\\+1P��Rچ/�B�h���n[����D�W�eWw�I�C�.jʧ����zY�8P��y�v�\���!҂b�c��j(�,sf��蛾k��!�l+�E�K������TMl�|%�ʬ,`��D�x�� ���1�(6�DK;�W�s���[�u�H^�EW����R(��rX�F�?^/�%(DǾH�W���� �z$�z���p�͙}�;��ƃ����-��f�n�f�P�M�JH��ߍa ~UH�y7r&&��4��\��|%w|�0VXm�#�H<���AF}/0]���e��6��鱼��?Wi��"m�@��U!���V����8�^:�(aIգQ�w��vBç�m�=CΌ��$�d����yLG����G3����k��X��h�to
z�8C����)(yO������+��y"�@�tW��s��_Y�g���s�SQ�LL@��DE�O�%l8��V�i{��_��*b�c1%��a�`7Ɓ�׾��΁tg(DH Τ�~�:~@*D>����V��J�m��S���D]��݀Ј��-� ̫.�)#:������g���i�}�;���P]4�����Ќ���K�����<�������-5a_"�s̸2��S�۸ag��[�d�#-�I�J��+7�}��.�)FZY�s��������@�g����Y�BF��Ao�_�rB��\�U�s[��Eט�����!m1L�TR!�Fon��]�h��h7F�p7rfZO8F^?ꨌgC~V�$���N\<����z�`��8#@-��₹�G�Ҡ��W�+���+^l		�	����%7|�$��۲R���Y�J�������pb�mB�Ѯ�[�&~.E7��?8�5��r�}X�J=~� *"�xUCɭ/ܜ���Fq!8�_��+��L�s%i� ���6hb3r]o�k��8��QT[�9Hr�~�`T�ņG�K�}���&�k����9��Q��]��!��o���*�MP��Ol�ۇ���]�sA^k�N��.�Ѝ���ZL��� �+I�Syo��!<�E�ş�s��z��<Q��'L�O9�]����Z&v~�U`м���s�[	�A?��WsOa��H唴���S�E��GJ:z.���E�&b�.�+be��f�A��I�`�O���by* ܜv[36U�=���M�M��5��Ć��m�+cp!����P* 9dL8���R��Œ�_�C���/S�}�
yq���TO+l��t�!�Ϳ,��>SN��ݙ�T��a��@�*#_-��F�!�DUVug�!�?H�Zy�P�x; ���}�9�g��eb#��]4>��p�;���\]�o���٣�¾&L��I�4��4~fv��;�
��n���5�"9./n��BM@���K\��H���;�+͸Һt��'�*�2�j��x�ޡv�9V��o�NiX��ܗ]k�7SVP<���2���嬯�Z��0P�)6k���R�f�<����yT:�D� ��	���Õ���
�Pal&���9x���b_������J&�e�ޔ3���P>��;�����k�� 8��W%2z�����uP���1 
]�I`�1��*ac3�%�E�#�Г/��)}f��HkD���GGd��)A ?��q���$6���V�-7�# A��ت�-��i�m��G�@g��M��e3%�[�ِ)�N�+]v"��MBn$�+w�5�q��񂬫���ܿ�f��X`*l�N�LпW�En�b�ސK���/���~J.�=P�1���7�C�r�\���D5aA����A~�ӫ�;�h�-�-��pd璸C�+�� W�ά���tu��ތA��j�ؒ8��t3�E�\&�J���0:k����5�%".�a����֤N�ډ/cIȀ�P��'x�+Q�dg�J(�Vi.=��XȜ��IP���Rٽ��Y����$��� �R{�~
��dP�qZݱ�(����\ҷҲ��h׸�����戥��1-�/Ȩ�f��^��Ȏh�����p01y}޼�\1�#
_�[t��/��&UH�����X���D��}��	���ar���'��}mO�1ܿ"�r=Ez$u�ˆ�`U���Mq,a�9����t��L�Y��V!j@���s�����dbD�ce�+F9[�ji ���[->����'�\�9��[��Ӗ|ݝ��~sK��L��%�d?5�U�T<�vj4u�`vZ�w�����Q����5�Sm�n��6��� S��y��)�� �X�c��gc�x5�M|��}#�w5g�OSH���l�O�(�	�r4%I����Ny��A�C�r"E�3��$�L�)�5�x������+*񨢇g|
g����u���H�<��$_O�?(�9oNy�!.���mJ�3i�T昗L�fv�K$z�&U)��(��Xkj&Q�Wt``p���1�.��(g� �<`Z�c�b"2���0u����GRxA�2������L��bb�K�����%��ɝ�쐍�ӚR�廍�)���Y�5��d?��+2����7!��ï[󧆄⨄�(l+t���F�)Ca�N���~��T���2[Ǹ���1T�u��͖%�Zѓ���ٵ��o|=�3��	)_Ij�2U�����p��Q�*�(�R=�_h磊N�j�K�;��ydX��c�^_�Z���ڤv��њ����HV_d����_�R?W7l0�u!��{֧�u�qC�f	�`�_Ʒm,��M��L�aF!o�JH� Hқ+U�j���|��Y�v ��v���G8�U�xH��z$�W��Ya����g&�U�lm�'�D�@$y�ѣL���n��`���Ĕ�����͡}�?�
/M�݁%t��.aʊ�쟦8�����'�Ο�d�f���P�n���g}0Z��Y}�����A7 M�m�0��;��O��r��/V�,V�=�h]m��wD���,̞���-OT3jB�vۘ�D�#��N���5D�MВ�Ԃ���
k~krJ��!^�:Y}�c���4-_V�[�B
P�a�Cb�TԬ�J&�����y:������N� IhGC�'L&�yC3\U���9Uʗ ���d�;l�|-�qE`V����X,�����נ�o�U5"�#��i����A����� �za�hH��i��_<wJ��?�qM߂��-�R��n�E P�8���h��t/+-֐��L�o��--ؗ�G��MF��	q2JC�R��_�Vm�O�凉�;���j�}B	��"R�`����7̆Ͼ0Un,���^'E:��E���p��J<�s�pM���0Y��ac1�����\	Q�^����r�����o�ZJ\xQk��=��_��>��Y����<�������Mh��]��}7-d�V���m��,��`X+����:c����C���䕰�l�U�{$Z�sb}*.�ZjFd]��"h��@f�w��Y�}`c 8�|���`��4�b��_�����ܹY�kYo?�}t�����S����{ �y���]��tl|�(v�0 3=3ݱ�oC�#L�hvߪ�1�)j~�ӧ1��.������?&/�n�T��!~�{C�����'��@w��5�t����Sj{Q����-��?����j��5�(~\~ϒ��T�u���(V9c�3Ц�W-� �T\��41����9�\��y�y4t����+�`9&�/����=�68vw}s�G�w����jS�w_,}�
�-h~�լ%	�C����2x���OrO�.�%}a�\~� ���R�_l(��*CM��&=�b�+Ǉ�����6nٴ����!�5��Y�+�����,1��p�$xr�9t�)���o&�;�������n8ݔA�g�O|��Kܕ���a��EQ��w����1M�����a�e!��3��|��[C�/��imlD���>��2��k�~�̻M�����d�zѩW�9� X�ֲ�U~��:Ռ�Qz���pe�X�e�h�ĂKd��"L��MiL��y�q�������X9;���~�)�튌[|jS[ �ba`�-��j��4��9���{���+V*�H��/Fz���F�ڿ̱����7zȰ"�Ii�c�?�,sZi���P��m�� �v���_Y�:LU[�o83�f��Q5�PLpTP7�@�q�ȨSU����6�R����4�_պ2vU����@ �_�종D��O7Я� ���܋@��N�#���ݥ�F��bL���>�f�F���*�X���W���X�n yЦKtR��2��J�y�jb"*F	YJ)ru�5���r�5��P��j��.r"
zLH�TYq��3U��T@:Mՠ�C��X�kť-p>�F�R��~�yg�'7�U��؄�|�/�+��Q�i��B���}{�&���6S&=���*��%�t��f�<)ק�#.Ǟ����GK��i��v�8��آq�]:,N2c����V��`�<�pnp}�u��Ňݳ
1�BT�L)snw�ќAE���C@�f߽�x�,���j�E�?�L�[��c�2p��7�I��"*\��`�5�P�4cX�dR�ɹ=���D{u\���1>�>�	V )3�J2X4�Q��wO��K�Ǘ�F;�P�bZ2:�׵���~/*�)W���nԺ��*W���5��F�8/[G��o�SVse���pG!~�zb�	*��@������n N=>��g|M�+6X�pS]V%���gIn�(0��� mg�m���bf�u$��
t[��(?e#�m4��>
�nG�^}��c�`�� ;�(���^H5/������y����=kY��E�hCE�-&�Г/O���w�$��m��M)z��*���;s����Nc�K��Hr�tA�1� ��<�@�����KF�"}�����R�������@<�xV�I&���k����|�f��̄��ydRFԝ2��;(���-��+��=l:�S��[���=ʈ����Mץ��)���K����"�U%�kz���K0R���Gw�	8��7����:uKC� <ڣ�J��u�y�YS�2���(�������z�5]l�6������ �ﰱB�T}�j����}�2�#f��A��{l	�D,�LP�эv�`��a�a�\ϡ{� [g3��DMSuc.���;����t���!/?I�3�i_�0!��	&]3��嵠���R��#����>����
ۥKo>(�;KuUH0)>���@*����:I��g��W7�ܜ�A����5���g��:q9�v��M�"�n���8�u�J>(���8+�����r��쭝��q�M5zr*�uleq!knD�Z(C�EPq��N*�* �HTR��=es� h"��L�>瑌��o��o|(GQ�$B��O�K�T�䚷����5��8E��)K�z2zf�~=�DU�<�Q"F��̵@$�	��-K�b�������9?�9;������7s�|�0�\.㚁���q�@T���;���SG��S>��/c'�T��27j��\Td�p���]�\�,�h���>
��8`Ǣ���y<��jbi��b�����^X��E�,R�v��̕�s��T���o6����m�VYcHoB}&-c dș�N
pu�ؑ޻ ��bka0XfW7�q'��	q�\^'u�sr�㪬����T���#��)�_`��-Og;��`P�2��s�\gSF����Э-�I��� ���M�Y�(��aw#��X�>4�Cwr�%u"���g-��r!]zj	��� �+�M`_�8�ƶ��e��3��#x21�X��[�QGij6C�mk�x�m>����;�#v-��H�K[��V`����Xп�m|��I��E+� ´�X����ۙ�?~Y~V/�F\��^a�,������;�\���a��#�<b]�#�N�j�R�.��u �����LX<���������j��Q�9��2@�4�B�v���%�I�q�%��Ql|���Ԝ�;�ׯ�>�+��Q'c�E��O�G��>j+#G[�[ھ��j����A���tN���R���>����=��~�Y����$ɯQ�Xf�Y���h�0`[�8l�Q�N��ɴ��# �d�'f��{��yq�x�m�Q�^� �����ڥr�8�.�o��C����Љ�ŨlD0�e�u������Ԥ<��CYNߦk__f7�@Pw��n�.Om���!�D
����̢h��w�m���S�5`	a�����A��9C��MԽ3��j��d�v��h!HS�e�Z!L)�^ʅK�|�|y �61�aR�����ݰD���1}D��ʵ_^��?�V{a|�r��a(�fl��K���5�	�:q�9c�#���C��	I,.������߮ ^s��̷/7�+���1y`��\��m���j����h��j��J���(�H���!`'sw�62O�?���r�z�����2����z�6�#���_�9�s}��ùl���T��������1Qzbs��T�{zNG)h�f����G�m�$l��;��cFxT:j�?pv
��Ԇ��1�Ψ���Q��Ć�,�)rV��*�j=��k��TNC|/"�
�_G��7:�	�����b�|����R�70e� �5��S�&~�n�ﭜP�'N8�yK?��W��F��ۿQ!�����;_�ǳ��9�%F[��xȰ/U��V��򆜪F�u�!��Q���rĬ�nEE��;��<\[��Qg��]E `5E����t�%��5헂��c�	���n�C��Q�i�qgGi/�Y!���8qr��!��W�r�_D!á�l�!Z�%8zRV����)S�#ٖ#C���n�s��dO hf;��?^]�̬�^�9X�G�u�A!�@ǃK�&U��ɉ9��rZ�h�K�8<Tx:J�[/�]�T��2������ U��A�k�Q$iq-;���Bch�wN[s�M�=k��$r^��-_�3���>�b���V��=���/��(�ajmz8����aP�9�DP[�n�xF�VO�x�"�C2�����(bL�U��Pɲ�n��
XuTh����h���YQ�*E���X'��7��U::�Ի�hN�ȋ6_�P�Tϴ����m�� m�D�@⻱5o�%���q1,уx���Q['�Z�zf[���s���/���]����ո�=� �v��0Bѹ��f��|xR��I�X|�d]�� �C�;�4����. |��5��v�$��b�:����N�M�m�m{�B+��Kҳ������% )��2-���޼N�żZq[�eT��)�M������=�ɓ���1��^EW��2�8�8�$J�����,�,�2�Tޝ"�eM����M1l���"�m`��A�&@��gc�u��X����)W�?v_��ƍ�˫q����u�%1R�-���v_Zu�:�V�דm�� D���zL��C�z[��)mRD]�����K	��˨�eu���3?OJ<���bDɳ�yW\�Eq�n���Y�J�96U,&ىh�]�ƨ��?���ΏB� .�V?t�$��]nJ�'�g�`�*]0#{ը[5`,��HAVg�JE9=j�5"�ζ��Ǉ���7����<��}�ȏ�����a8q2�	�g�F{���VA����֡���iO��f~'��wZ��Q{5[u��"����3u��jb�l�Ϻ��.sr1e� �)3�9��M#�܇ ݊�+�[�ö� �A �V
\�C0W���6=�E�&p�C.��͞Hn#��+R��R���~
��EL6X�f|�Ϣ�tM���o���|"����C@׻��O�I���=�5L��ڔ�E���^>�;[�x���K�����?��p�y�nf08��*\���YM5ѦRs��9� �>B��� �An)}���Wh�
�W�Lˎ|5.���>ف�WY�a�&0�
s�|H�hY�z/���3�i�y!Q��ߍ�d�u��x���o iE�q岒�ӧ t�XA���A �䧛�H��(��)���@���p��s�}�ϳ0�1a�.���"��e�PV��Ά����'&ßR�Ty����su�`Z#�m�z��B�j�����?���������IXT��QcE�!�7��)8g}�&�Z�R�+i.�Ʃٸo�h�&�8&��A��V
N�t�ʹ�G:L��������.V�-}t��fk�=c��ۿd"!"���X7z�