��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6� '�7mF��+�Q~y�[?(rЄ[��H�{���Zh�ƯD	C�o��M��+�I�J��]<At/E�8~�8Vp�Ef�'�ǫ��ZW� 	�,�*�Y�S�gF��ӏ��L�2��-�ű�p5.Ha���H�1���� ��h�ڗ�h�|7�F~�QNy���RŻuC��m�4#}�ND 4S1H ���J����Ě�XaȚ��.�}x�M�W�[�w�	Y7�65�Y��6�4S�D�c��sA��!�Z����BJFAϛGw���V~er��k#!�19'�^G��N8�9d�~U���3����R�be����w=�O�>�[��n��U=��Z_M�@�:%�� �y�{����he�������,}Z�a؈�_�y����e�I0"uz�<�`v�2�Ih�����aY�q��G��4U®�7���u�Ya�X���SLX�2ո�ol��Iٟ.�zSoF:,��۟3���Kq{���`��Zȡ`U��㊿M���o?6�ɍ�wp��q����f���������o|LI�E��L�(q8%8�ɦw8�aՃ��ÑP�Q���Rh5̒ �AP����P!�R%5�
�^d����T�#��$�/��##ݷ:6�=��+��[[i�ڕ-����oXc,����	Ѝ~��"�'t��G.`���Ru�_�I%��܎<��;�?(���:�>��de�3���w��E��hg�\�D����M�g;��ϛ��OC��B�ÉNj�ƾZ	k{��7�BY|{?&��{N��GH+�};�)撋�]��N�p7!�&��
�w\Mڟ���D���Q�`���ʽ*R����=�<���`E f.�6֕��]�e
Y>x�a�Je/{��Ó񗄹c��L#�n���kԪ��%��6��A�x������11� ��'�?-h���N�B�hx�d�z�ؗ���EE�k*��"�KvV�b�3�����c7��U�Ӑb�F���İ�[T�c��)����)�F��wr����BH>(W��iZ���g�~��1� �X�%G������D����o���ң�&�s��[ ����������,Eg��^�$�'ù��V�~�?���3��S<C�0��~י�Hۛv[�r�ïcI+�;W��Ѕӂ;�?m0@
����ܯy&�L�xE��y�G|:���ְ��#D8N��|/�펾V��BQ����-
V�!_y`�
��JC�X�6��紸����r��wE@���.�:��(�~�^�>a�Q���^�Qm�
�y�{�潬�����*�{��A}�g%�����"��z�R�a�e ��w�ص��>��U�l���Ǳ�6��V�˜x39hO�B񰉅6�y�P�p��hW��Dv��2hh��M>1��26GH��w��,�)w����Dًt�����zy�~V˚`��R'�e�:)CF�}�T#Ro�F�����H]G�p�F(]!d}ߋ�a�m��ԟBȰ\�0.%ӓ/������t]�0>|	�8w��du0�4���h���1��)S��7��0�4i�us�/9A����跞�7�W�E�#�u��g�%k������ک u�ٛ����~�S*����k}�-&h������*������dO<��l���]�5�KzzEH�L"�ҧ�OtOoP����a$W�8zwxkH)�J���7쵛�����c��c����rC$j v������{��{���M��"n{��L��C�ʍy��ͽ�b_��?܀ٕy�*$�E�5ՓP}�����T��	M��Fi��t�`J�}�\5;�z��Y3���4�f�P"'�qx`�g������#�=o|���t�ߥ.�/8V
9��L�yK��U�.xB+ߦS#�E��y�"(T*��-���&,<H�!!��C������5J\��9?&�d�"I�>R��ޚ�2�K�E:9c��Lo,�w�!_�����t�c��G��M4���m����̾WYiX�h��I�_9����I��r�K�My��jЊ�MR��N=|�	�n2ي���J,�4����Wm��C�_��2�- kj ���V�&M,�K��nQ�ʐ��8�Ed,"�y[����d�����TѶ\���������ӅM������[u���8��8��X;�n4�`�'��D��������ia�+:��,6q�'��_�vלlr9[���/�a�֪{Ny�z�6� ��녒ld9�j�1�2�=(f��Ŀ/y��-ѭU2'qC@��!�Q��!����'�����d!�b�%?z�$p�����g[��W��axܕgCD�-�v1�gT,���X�˒�Q(�� L
Y(��z{��D����ΰ���sԻ�p�ϸ���-��^ܜ����7�lmI��
�$#Y��p�g���W=��4N������y�����:WH�Xz@���ܒ:�����������M�;)K�b�fn/��^�� �p L�iwj�HFhnl��"�!u $�����_�����ʉb���+U�:�鮍���۱QA��d��>����t���z��J�� ���z�1c�(R��F��!?�� ��3�8���_o?<�,JсQ,h�f��?��IF0�Q"KwX�Y�<P��Q�gO:Wx[Z3�R��t�p(��ox�P���� _'y�q.Q��OH=b��]O\��*ĭ@��uK�4g'��9�98KXd1�>�=-����*m[�Q3F�.���c��A���
�~#�͙ ��oc��H�>PzW0�:����N�Z�BO�9�T�iگ�WV7�?G�C}��VM&]��R��e7ȷdx�4ޏ��P�$R�G�wmaS��kN�[�J�t�fV1�h��x.�/�����ϵ?=O|(	�=�� 	��{D�*�~��,����>gІ`��
d�a��0W�6�pG7����z޻c�r�wb�n�����r����:�ؕ�h@��G�A� ��*�S�3b��	0��2��<��q�5��&�t�Ű3�H}����!Ze�ȡ�s�O�����>>L�O��|G?��dê@�S }��	��]�e>N9\8��i$s�Y&L�[�%O�s�<Y��SH�Ft��L���s����q�k)3���G�����g���2�)u�e%l ��?���䏺�H߀U=�*����(
<�R�F�LV�����$po��1%st3��t�m��%�,n��ڠܬ�ɭ*h4o�����/3�y�NeX���zD�	��ړԾ�g	(��Çq�f��}p4�)3�g�q. 	U� ��J�唀u����Ǧ����jV���U\�Q�R$ݿeY|��NX�� iZE$���Iz|�Y6n�
��$� ���^�W���PZ5����{�	���[4���Q��>�w�U�NNLxAQ KZ�&=�J,��(��4��Xn\S��Z���Vy�2L+�Qܫ�%g?�;��g�;�˧֫�?��"x��Z��8��բ����E���&k��U�H."�;/$�{hϏ�D��t U�%�`��Z��Ⱦ�<y��C�4�#������L�{{-x)_#EkkҢH!	�c��n!�̎�VD�e�!>�y��l�����3�[k�P��d�F�@'G��h.�6���p��%��I�>1�J�p^z��eW$C�&w>:?oo)��>s,V���G�6��
�x����Ĭ�|�+�u��,.�c����г���#lw�v��Vj
UdY>�o	g����N@CBd��Z�uSv�]�����qЋɏ1a�g�*�)XG6���/�j{.&���B�-,�5U���g˱�	�c�ǑA�i���E���TT���C̱���ƺ4��U�A0�c;��ʷ�@CO�=�����Nrw�'!_��U ���ȷ������X�j+�m_ҳ)d��E��J��1�6R�*A��Qr3	�O�g�eK������s��@q:U��.o<`� ���r�~�:���Jo{<�t0�?���X�v@�R0b�Gp(&�­����K��=&��?%q{|�y����O�>�N����m�������Y��Ţg��Q��0#�^E�k�	��nLmJhg;��jM�\Y�]J��N��q��,�(���]m�P��'���nr��i��Lc.���tI�cf1��Je�/�����(�L���I�h�?݃,h�a����o��8��i�.,o�p�J�\[�pA�q��v��"*w�cb�'���������?�'P���i*6�nwz�?��z����fR���*ĿLHp#�F��ԃpf���'���#��i%�B��3)d�ң:�0<;P,�	
[y�_Ĉ�V��f_�߻�r��K~�����?������ ����SP�t�{�K���'H<Z�|?I��/�c�%�+��I	���q��Jdc����ٺ������e���oP,��_Ihaɨ>1W��?k)��&���N�\|H5�q�������;��
�K��_�x�^�/gŻ�
_����1��Y��_xit��ȥ踢#ݮ_(�l,0b��n�bG�L���/�e��Ӗ�<BB�]a�b(�aǮ#��q.�mׅ��/uC6�����Z�V�����Z�gtgM���l�E5|�����F:��ժ�s!u�eZ�!�}�����aM6�o�ن}q��R��
}HQ�<g�&�)��yÁ2�on�v6�{���d/��b=���d�]1"��Z 3`��|T�(d���r��u��33�?����� oz����3P��7+�U��|o|&�S�d�M��s�S ����Cc�hq�Q���?�x����EM]���{|�7�=�����%YNjq������c񰺈B�\4Րw����%����`L~�y�������?��ʦ�S��)T��u?$�c"i�t �|�߸*��Y��B�k�����:�tE]��I����E��橿��Y!cS�D� v��o� �4�CY�?C;#������ּ����q>��I��q���U��?ֺ�?&w��v���R��d{��h��{�o��;�'�}�|�C��.ق7�#��0����&tyf=����[����f��ۗ�]a/��H��;8&t�HVWOj/��ǇAE,n[�ko2P5��K��-g{�B ��󟝬8�J� �mz�3��\�0z[.��{�Ðq!�>*��W%I���*o3㔋�4���eW_�qH0�6�v1���d�t�`-l�d�؛�jli�>l�7��Vպ^Բ���
�l��1��'�1��B euB\��׌-a'��6�8(�R_�������P���"@r_�C5x�db�z?NY�i,@$���`�Wۖ�[�IyĐ &�'��#�}�	U�S3����Ek�,c���ڱ7󠕀��$�N�|��� FZ#m|
�D��J���aׇ�8��Q��k"�#���������N��!�A4m��_txr�?'��hB��3ǲ�u4���zrL�a�:s��෰��f���kQ�?�j�>Z\+ob+;�����I�T)@Q�x�y�wT��P� 4�a��!�#E�1V���e`,'S��I�
�x���"����+M���Y�4��n
^�Oj\��vF��t��]�����aJ��[+$�o%!L�ۙ2`U���k���T��?�Gԭ��jh~�N�+$y8�B./W�,3���?�K尀}M���MW�mE.>]&W�D��F��4P���'%9�b����t�o�p�������3�ƨ�]bQ���M����2˭���G|��J9��B��E�8P��R)��cM�إ��ޙ>YƘP(�:D�{Y_���~&.Xx�8��Y<��IsK$�V�i������r!�}a��q�0��왡��9�n�'�t�~^����C' oU�眙�T�	��:����"^<�+��P��Hx�V3�,�
��������M���Q�	U��O����
�So��� !�SK1p�����h&fxNX�_�y�#�?j�V��+��'�t_~Yj��b��g��j�غ�d&]X\S�7����\�ޫ��O���7qJ�п�,�"O��σ�k�̖�\`0/E4�k,�&�x�T�)͋��h6�C����TEV�(���/�f �u53��Aģ���{k���Y��`�r��'��K��3������b�����	�1�0�u��n��z�2��h����X�^V�U�y9L�̦�ZL����r,��yOY���lrO(l>?�<�&��w$�}
��2S��?xݜ�Ib��1���
).�b��<O�é��	=i�s��%e�����ݥ,�C�o|֔��,{E$�t�|�x�*���.dl����EF{>4�%���Vp�,ka��0�=�c-�16W�]��#������-d�;����O��=���;o�WO5���:�x� 6��]�y�ׄ���r��n�!f�
��oC�;Z�CE��h��uM,�?}�qt�0���k�Ր���А��A�|��=�q���K[.i67Mpgs�~�_�E�ֿT$n���)����L�O��w+4(�8��Lfyɘ6\��I]����4��G>.�f�쮘��܋p�x�j��}����K��݈��Š���v^�C��<3�C��u�KSf�Mqg�tLn�}̄����c
�{�'�i�$%U��	A�
�3�kM)�ݧ�08 
ba#��TZ�rզ�J�p�e%C�fIY��W����,�����]^jੴ��DW�#�IhT3o�3�v�ZYv�9�d�#�y~g������m9cpỲ�J�p���a��(�;�������阮T��]�W-���e��}�q�׻V3�7��UR���S�g�-���۲��j�%c5<������ԭ9�:�M�*���0s*m������Z#E�/������}��xl?Ih�4t��3�bZk̕B|��>sd�K�n�T�v�jٷ�Y����+���A6%�і �M�4�:lmlgC酮�T���؇�K2�v���C�l�����0v�s�nH��GRT��d0#���mֺ��	$�*8��~��
����T�9����}�����8��#�V��R�z ���-ְ�;!�p��j�ɮ$��/�"��;�H�슼%�7h`3��q�_'vh,7�o�03\+t�6-��//|���%Y��皒���.��Qd�0/���1;��IC�d^��)J"c旄(b��ܒ�OnG(��o��Y��Ȼ1��� h��ܑ1�g���_�R�(�������4$\�u򈝠�)���i�u������nq���"���P$��Ș�6��=�`Z����"�NjԢs�`e���f4�Ҷ�D�^Z�R�C93�
����S�vx�!����� ���̥/���s�cEQfj��.���Z즐�_����JV}��QJ�p)����g�����;j�s>�H	����.�O���Z�s��z��=��j��Cv�����<���e��Ġ�|£��/�7*YJeǜmŶ��I\w�OΕ�fd!�C���N���MŸ�w���d���"��|&ٿ��k^ǜ���G\43 �k-Ky�i���@@�"{���mbX'���i��m�]l(�ѦfU��3�}�S鞗"u������T)5�!��h����Gf�=h�|n��=��U�7�P{�vsb�>� ,����C�~������a�tV����=]�]��@)�I;f������!���aw|S'�[��T�Y��J�Q�"&��@˵�9'���xog?)k��gf�$�~��<�5���G��D��gz^�za�0E�m|����Uٌt/W㩒��]�c���'ߘ�� dL��u�l���|��x�+4���F���f&=�@�*x&��j �{b��i	�qf�9uR�����T������������.���\T\�Jg-h�Y��DB$:I�r!7#�걯1��`��%UZT��qjN�x���]1�ͦ+��f�W�7n^�z�x����`��{5��'<h�4������1��	�]3f�ET�C�ԛ�Ą�%[�0f��®�=��f=y���:�f8�R�ɸ�����̷��D��]�`�w��s��:=].�uy	\��;�$l_1�%��Y�	/u��eʳ(L��*-��Ջ��!�d�@l�	�F\2���"� ���`D8t��^C%݄�V�\�$�=�wvTsF�c�SR�-�
�x~���(��Q(+�%[�R���v�Gʤ��(EO��n����+�O��G��&�Tb�s��	(f�����g��#F�Fe7�N6��)kڜן ��mT'�ݑ�������� �40V��!C��
q2M�ޗ2O&��D_!Ƽ�#-�r`*؀Bwa'�>K�O��$D���<e?8�����y|PyỢe6K�g�5������Y�	b�K��C�ejk���V�V�@��ۋ������;�J�����aP�#%_�gp�-�i�c�n�ç��H孚<~eR�h��;l��1�z3�i�B�`_:���E¥��W�gG��]��,�x�(d����3f�s����h���U�]��Vq���;(��?�*Od�Ol�,��kCFz�ȿ.�F�>�o]
��N��?����r�>$�wB��f%�_ [Bs�0p�b&bQ4�I���hV&�ψ�:/��6l��>�s7~�"l�mX��g��:,	��'a��˴�2�-L^uC�3��l��`�E���/K�R6�}*��+��H8���8&,��%B�`�smϷ
�`�~ԻLݮ%�h�g�5$a��Č4,܄WQ_i���lϦ��0��AG�<r|f�F�6����H�
G[?*{��Ѩ��{.�����.F%&�9v\���bc���KIB;�}�Kt9��l>�Np�ut��w�6��u�l�!˥+��U*JH���~����"��CFЂ�u�i/�}@|�J�ېǽ`W�pD�R	��A��Z�PS���IE��I�k�Q�=�ς�#�l�#L���z$[���،����̅rL\�d�JS)�e��Z{�� �7��Mꠚ�M�����]Lt 8�yK$�"��RbNycV�41(�	hF	L	Of�Uʳ����+0]C��ޠ���,��{I�#d���۳�=�_�
uKg	��h!��7����70�j�C�q��J�nb�J�MCRە��:-7�Aՙ`�ö�Yt�a�Dt��G Y���.b�nLʒj}*�����UJ����:�����8L�~�eI�VpD1�rN�F�F=��,��+q�!\��~�*��|�8�aħT�Po
h�&Ȩ&��VFu"�w�LM�Ԋ�ќ�A�f���<�_ΪAs-�k�<�d�ghֳ\�P�(�t\�8�[���l����A$��nJ��1VV��(:&dSr+��5gw4^��Fk�A
kx̨�r��I�(jP�l�g8#Y��fd��s�����G�R�ŀ��O%���@}d$�^#�zc���RR�=�sL'��6�$��mQ�-�u �3�kK��b�x����-9�2���kQ��@T7.����0%l��|�z�҃�J3x�`<�g]o���(��C�k�_���{�`�3�m�SOPE�|�=��Q�
��A�b!��\�0�����p���5~�V�����o�K3�1'�٫FSS_�<�O^~欮pȾ��&����F�`9��"O�G�����*�@�x�*0!q�>ץA�gs���A�<m�>A(�A}VM��_���*���ʈ0�9M�ua'E����r���%-O���+�����Ab͍OɃn�kKW ��e�<�!<˩�j�g���F��簏������� ��er���#�f;b����kK�N`���h�H�fvz2� �1�Eʦu��U7��f��FB����t���(�O����K[)�k\Wpܡu�@U~�S �đ�W�X"��0��]D~;�����h�]|s��
]�f((�4|>��	ʚ	&�]q��qjl�a�������!#�)�<A���Z$�����~�51��ЭL��09����$��Ԕ)KC�?����'}��
�#C>�=�ެ�/�Y���B\��,��'��3�n
��݅����+}����.��$�}���l=��2)]z�g�}�����@9���<^��I�};��$9��N�h0��@��P��,�?X^F�fG8ayW�(�X8�NYP��G9�翷
7Sx7��Wk�u��2�H=�H��+���[o�!d��+hඵ�V�2��E����������kE\`M�a�biu3t>���c�Y:*p|�J�A��.fF����4Jr���K�#� �9�_�c'p�LY�R�g�������UC3
Xk�N+�Yyg��(��q���x7��WXȏ�L� |�2£[���Bؐ�<^��<34(Ѩ&��� ��;;�x+�װ��;��f�����
���������o s�+X�DY'����h�Mj���hF2N	#�<g��fVb�EDw�b�)R�[[�P|u�@����r.�#�[
n���"�2K(���]�LF�Tn��䈕���5T��∶E[J5���K�m�	�w+ani&*G��b�=gfN(���$�8�Dg݂~YR6O
	ץ9(9��FZk̈qhn��o���|�%��˷��*N�y{	0s	�5@�L��!j��J?���"w��Gc�X�o�c�8��6���~L�6�Z���� 
�m"1ɡ��ϮO��>K�x����m��rչ7Yu��m�*n+��s*����i>����+� ��d0��B���(��N|�u5�^�JQ]W��W�k�F����������֟lf���2�85E\Յ�5Q��D�7t���2�{d�\X|�^�`�U�f�/��g�����A*�1E;�H���V���1�UPi;F5/��?���#A��K�'-b�ߦ���5=+B���="�QC>�$DP��y"����[Ql��~}v�$&o�	���\���D�ơ�'���u���*�d ���r?�(�iLq�h����1D���=n�;�|�/>����&{�
�eV�䧍�1e% /:.����ˈ?P	��Xz��
��S����/>u�u*�ޤI�e���0N)a.����Yw�l���Gɉ4�r�c�|��_��ȅ���rEA��
.p|H���e������P9�F���n��F`���\\ \��W[������*tPx�/����㹿zgON���A. )��|��<@#0qZ��=��&���P��Z��?51���;{��
Ў��f<Хŕ:�OLܠ�I���<_̺4t���|ϻ�%��}���Pe}�9�z`��"�,��]�3.�h�.t5z�ʺ��nk����b���7�*�s������dZ�H�4�;�ZL�7n&,�-8\��@�E><�[|![�_Kj�m!����c�K �F2����:TX~ؖ�D���b��)�B'�`z�&Q�RcOj��-��ٽ�d���VW2�k��݊4�pgF���X�d�;%Z��'͐����V�+Z>HrE��hhc�`	�;B#���I<o���F��,A�ف���@��HYh,#��#�.se���N��s�>����GdӮ��85Zw�o7����x�5����)�O�+wFDC�6��uU�f�e� 
��Ip��(�����	�EK2X��aE ��+��~�u��݀n]��Amh��M�§,K��?��N^L��J�S���N7�B�m�G�L;�Q�l2��?�S��i�2�8�:�[8|�y��o�i���}��J`Lֺ��� ���Ǟt���;q����m)�JF�gC �Zz��)��إ����S�����1��X8�9`�H�r�i�%�ִ����Êi����'a�wmq�H�����~ƹd�5��B6�Ws��oR,E�Xo�R3�T��t�,42���XD,t�4�����Uh M�U�BG
MP��:�`��a�f;9T),�y�W�z��pZ#�jOT����ʢ�o��A��p�;�5��^$=�?�����1!2�N�]h(�oUŘ�ܦʓFT�������+v�m�ˍ�9^$?ip�L�s`�wC�A�P�va�U�9t�V-��ġ��1PĄ"bˆ&�fU�X*Z�Ѓg�0�Ȃ�����*GUD�hK�B�N�ʎM�(�$��jD'���G:������ſ]e���3�y0������t�<���x
�-����ruٕb�0�2�bB�ߕ趀���u�/A�\�ڲ�S����L
_����9>,l!�0���۬�"x�mY�e_r��Y�h��S��c�q��x�܉l�ACm��n���  y�� g��eӿ�#I�ߩ��k�0 �+�H�_��.l�.�e��P
z�7�73K5�sw&!�U1��6���k�!�W���Fa*`N�O���<,�SV�����������(�{M'tyc��2ڨ*1�8L	�	GO�E��5}�>9�W�^4}��:����:pn��sk
}x$�9Y�b{�)G�R��w޾;r��JGU����z����
�A�$Ӹ��&���rh�`��82񲙢����1���;.�{��;,u= J�z3�n&���YnBڜ�d��&j�}M69���{��T�L�~�aWc��Ј�E�Z�O�ǂ�s��_o
�Zw��-�Y�yZe>�^�b�h$���w�o���- �;�m��sw�hv��E�~�F8r�w. n<�;��r�E[)h#GӟO�@22���?�I=T���g<W���H{&���x���]"�z��CO2�����!�y
Γ�:)$�T�y1����,�>^��ɍ�T��� -�$w;\���+���p,e	����z�/7.FYU�ȧ���p���ᘵ��s h5�,�?����o_N��Y��O��N���op���z�}��%���)��B�`v����f�;=�M��W�����V���yߌ��ʉpX�"�4+V��l�[R�=� t�S�}�`)�����{�E�d�v+��	�=��������~�2��"es��'2��?�����!�4�o�Gγ��:�5S��i���q_*���~3�1�.��(#v��I�U.��#vIU��;![8&տ�8�7�6l�i@`����{����4���k�.rW�%�w�o^�a��X9��;8@�-��\,�ؔ'�'���*v�a >ϡ�5��N��_����fr��M8�ȚF���YͷO2��`�SA������L.��W:�n�P����E���h�����pK�ǙЁ%u���W5�����N���܉'� �B�$�|��� 	XP���$�lQ�8�9k��mPC�^ߖ�D�
�4��+�sXL:)O���n�6,Of�y��ŁД7���J���RHVg}Æu�thJ�U�ʕ����ʹ�R�f���s�M��4��?30��|h���7Ǔ�|��r�8�Q2�OgZ8���9��yp�c�q*|��w�>�W���]����]��VJ�X����M�����K�����h�q�&�=�
�����sΜ�'7�#p�Z���Q�P�v��*�Zk-�n�
�������v�ȥ_#�",á@�oP
�JR��T:� &@���+4���'��H�����-g,���L�~W��4�o���Eȵw�;����O::S����U����Hl�x3����[f��3	Z���n=����w��1v?��͗Y5�)�QΙt�ѹ�t�&����ɨk�w��K�־��0�$�hH���0�
8aUh�q=Y�O w�F9�\�>�^����*5��+n���V'>�tC��i��g�y(0�HS�i �!�wH�M���{����,H;��=�u���g4Y�EpK�RYҮ�Ⱦ���*<LZ�^V�X��/���#Ip�*k��o��AJ�N��ރiAtZ#On�m����ߛ�.)N�)� ���c��@�vr5+��i��L�i!�	�6�n����eU��Y]���ά-`.©x�J3�����ǰ7y�'�̔���en�P@���0��(���ٴnx�m5B�p�Q���x)r�~(���cB	>o�U��ZF�2�q�4�`u����M�{V���]�L5L�&J�yW��ŅN(|������� �EC���X:�H�ؽ_N� ��5A�5����aޑy��8骪N�]�z���tq�[����	����hsi����ܴ
����jLu�]�*�LSK�2v�N��s=T��F���sZ��ipT�ofdj��F�yGR%���5�>M-�������X�|�r��%�!_%�z*��	�|x�at-[��r�(r*͘G��B �NRF�m�_��6�R�ߔ�7"8b*�c�0?Y�G���2¯ ���+�ٍ�����b|a�m�oG��xm4MU��%慥�HT]<���X���ʐ*p�)'ϫ�39���E0��R&=���(����)��+�f���xZ�����|�ӡ�{��7C�+2%Ӥ������[�pe���6�r�9%�k��z�AUq�S,�l�@_ڟ9dXK����1��ʑV�$�5ھ��`K#�|;�z��U��2�cߝ<_���9"�?�è5e�͞��ø�]��� Ks8��6��M��[��iߙl�J�WN��j�}[:u���?�W�_c���˥/��=�˱b�ft�y)�^�H�h�6�K�>a��0R׳$��,�(Eڞ�aM�zx���^c�$HN�Z,y�¦"�xs����)�;�[���׬��AC��J�K2f�\9(D��y(�S^Zb>_r�",bL.���j}ˏ����y<C��T�ўh�F��j̍}0M-gŐ*�[�SZ�V��_J�����<��'�o'5P�4��0HK�$h�-��k\֩�st�fkz:���J7�>V� B�0]@��mYS��5d��ث`O�S9�"��������1_�|�9��P�iI�h�Ap.p� <_�"<�r]�-�����"��'}���Q�f�_t�!������0���D�F2}dyJ̄
�xO(s��beU4\��'0�C\o-3&��g�d�R�_�F����G�]�|Q�dCs�k�Lo<��h}���={ ���ⅿt������ٔ
;��#iЗ���dr�ma�c�:z0CKX�de	����)%t���\�w�XhavI0"�3�ߞn�@�3;�YM�̽4=�:���y6+��ՠ�F��X;x��aZԅ�u{a{"`�|��ث6_��f �	�'���?�]�y��^!���J?/�	���/�8�[,p���U[��E
r0�SO݄���t�]�K���D�P#S6��Y�Ձ�vBރ��Ki*��M~��
���M����7Ba(3���v?�~E����~���[�B �*b��X�o1}�����vpy�ϋGN籉���Dۊ)�f���aq����Ci���ƀ �-k#*�҈�߬GKW�9/���h-GpX'X\�~_do��q�	L-�~j��g��F�s�K�ET��d��ey^H"v����������yb U��}�Jc�&zh�g��������S��A�%}���`���9P�7~�J�rt��<��{�:P�Ml�*�q<mr�#N�B-gϑ�����	�W�E����Cmv���[a�o5Cv����}�~4��)��^�#�{�!� ����q���N���ʾ�g��({�K�rg���)R5i�+E>2��t��]>zM{�c-�A �����><��mz�a��.��5���N�	��ʑ��%,�O�{5�w�9i�?�~���Vr-�?Jus�Y/V�xZK'�%v��~�4!`�}�ߤ� �
+Q2C}��v��;dc�	P�"d,���~
�c ���yG�$�+g� ��|(b)��J߰<X�ϖ��u���O��0�4��Q� ��:RrvNP���-�/����,�w�C�hd�S�K%6#Пs��Z�8Ǘ�?Aq4J8��:�\�׸�:�rǋ���<-%־�����!��i����pi���v#�x����v���S��5�+~  !\���Rя'�z".����.FagN;�gF-��Y���Y#�8)���)M��+"�H���?A2&��7C���W=�$��ߴ3.X���4/%ϊc*������j�GUQYr^R����G����ģi�;�
@p�Ɲ�G�1��%$���YPn8BBMn(�,VMJ5KH%�-h�ܝ�kQ+K.��1��)q����]���w���G�*�����UF	�+/"L�i�jc-�9�Eޏ�9O���^�1.#�l0�H��1A�`WtgL./��c�����F����-è�K����f�xR���z�_(�Ţ_��Ň�	�@��?\(���>Y��K%��\
�IHe��dxn�7�1K���̑��MU�a�WBf)XbA8����������b����;)���?j���=�WB��0�a:fS�6Z�{:�z���B����"���)�����<���+=����F1/)�?5&}.~�����qa"�ݷ|t}X�]K�}��j^�ϙ��}�?ȸ}i��Rxu7���g�+�AQ���A񥩽$���
��q6D��s5��Ȳ�U?@s=j�Ӯ�Y�Wq��Bep�ᮬ�1ӑg?;���Pؒ�fZp�b��c�'SYz�?�d�@��X�D滨׸r�T�[?M*�!B�Y�]01�珹b�BU��&!��xxO�Do5�R]�X�&J���.dPͲ���YxÉ.p�Էw�����V��c�^�e�2j��!O�܅���B�k�dں��L9���ޖ��o$ءQw�q����	�鷴}�.��y-�q�ϕ-��0��?b:F�2��-�r��y~)�_��������>9Z'H�q��`K��l�09q��c���Je�oV�����V����y&��e�?��]O��眦�lT�®?��_�M	S�ϕq9�׫��Έp�E�`6�L�?Vc�AKC2e@%�\�Ls�§[?�;+�8�a�uj�a(�Kq��=���� �`Z���I@[{�� �(6b6I��M#-ד��I�˙]}����)򣙃���SU����]hm�϶@�aЅa�ڧ�p������K�?T�b�I�	�u�OT�~�)��9���9�ߞ�X��xɝ<�'�\%:�����V�bs�E�J�gU�+2��WU9�$eI^�x8�q�Ҍ"�͇-Ea�1&��NO�n=����M<!_���x$'�
p��(��5Jzg��t���"y��}]�#��:|B-���6��R�ZCm�P��,ͰƏ��5�k�ָ�R�4q�)G��˚%�l��;��"�(M�*�>b�UrMKxc,F0,�Tʗ[�Qq��Pv�E�m���]BU��4�S%ֈa���tq�&cHo�*�������2�~���f������Ą��5�?z�k�&ݯ|�	8y�� d��=���GDpx�8C�����ay_�z1����'/��:�;ӻ����hF������[8{�<h��{pE}c��ӈ����+�D�k�M�,�vS%���a"Z�ր����Y�f�h��c�>D9�4�i�=�6ٺ�j���Âin�{��E`}���

'T�l��@�ݢ�[5���p�*��Ч�Ns����������{"ԥ��:T�K̙bs�]&���E��X�~��?CJ�[��⥣۹��J}ږ5�T���N'	j��E:P>���M���]��zr�U��-�m7��;B�!"�㩮�I;���}�vUݎ̷8BX�ȡ'�0u�/�z�>��E���ԫ�Ơ���MyZ,�`���i��3خ��el����`�ԍ�w��f�|x��V�͐c3�)��G�h:�������)���_k�[a�F�Mj�',F�2N-���Z���у������ZҐI:�Q��*U6�(�Sx�8�5��p��Qha��!��x�B�5�ϗ�K�(]D�;��ebPi���=��g����΋�6��c�q��1�P����Uh�A)�IY2n��>w�L�j�y����'����@���p�k���f���GU^k}����K�I�j~��ήDY��G��!MF�J+_Fǆ��x<CY� ��J_� � ��K�ż�z\���D
��a�����i+�?�P��A�^��z��V�����){dh��o�9V{Z�{�_���9��Aj��@�,�3���>+B�	G��l��:���_~~�G�F]�#�$�'w��`}�:q�b�H?Ä_��!��\{�q��r�R:��
��4�=w� ����r����rc�}��-���[Q��}�����b��}�0��'�cA����@ܩ8ڢ~�������h�5&�R"������#O��Q��0\,K�Ι���P�С��.W�I���8?R.��9�Q�նt(�o�.�i�1�@4,�Ek�Jd{�k�Y޹|7�)b�1�Nl���ξj:g J����%V��������Y{/U�����B��D5���-�`��􉇛�9Bm�!����N�Y�WJ�Fo������#�P#�apqܴ�M�Q����R�4��b'�į
��K�a��㥮Be��e���Q�s�9�N覛�p&�9�A��6Ode3�s��z�p��5v�:�)�Sԃ�xm٨;�8�oM�-@c�)���r��쐞>=��R��]���� �\�҅��$��L�'�͇�[ӱ��%�84gk�J�%�ރ�9$*}���Ȁ���һt�P��3A���^���pԜ��0]�.���b�:L�.-U�/EQ	�N���G [���y���x���� ��c����]�ظO"!9yH�|�3PGxz�0N��iA,�3H��=W�w�(ӾY���'ܚ�=A�T�tR�LT���Ǿ�@��rO�j���Tmzͪ#�V8���ƫ��2��v3=-�lo���WM���<s��S[�M1�w�=m:Ϸj�G4�'�V��6K ��b'���Ѱ0�}/�Q�<���,�s���:K��
(��=E�����=_lrg^�_���Aѕ�p<���m��0=7h��F�G�N��!3�rx�3)� ���V�P\��#�<�pL�^��q�6���Ƕ�U]I���~,�#EK�F.�[6�.�t��=m#��\$�����; &��/s~	E��q3� E��J�z���i�l�����)�/P��ָÜ*��x&�<��D=f�SR�j~2y�v�3~[p���{+˩�~p%��5X$��*��W��iɹ���A�>$O��H�3=���?�Z���w���i]NY���iC_�nH��j�l�$8V$�l�({4�D�AD��j���C���i#Vy��P���'g)[���J���
��"%T [�Q����@�HdY�Rm�`dbK��o��*6�:i�%�\��p����}�}H���@YD.i��-���6���ovh��v�B��q_��1�"��eI!+�kA����0�QShi�g�7X� �G���$<,,���o-J�
��O�����$CR����|�lBNE�]�T]�I��q/��
���2DE��Vx΄�Ҭh�Þ��e����eC�b��K�v| �ז��ܮI�=i%K�5tbe.��a�Y1�"u��[l� >��E�Bc>2����kX����昣S��L�|�B�*�)L'[I0�"�ӣ�خۋ�#1Ci$�9�c�sT$'��*r�&����oh�%��k6�9��г���c��,�_Fg�&aT�ydA� �s��씘�?.�,Z�O6� �u�N號M��׼� &Ykp�y�)�X�y�v��֏��Z��f��L�`3�$��-�_�^OB�s����5�*���[�2�JU��!�Ȓ&X?s�+���-,$����k�5,�Q�z�l2�Qԭ�M�����DPq<��7�D���n�,�p��-���S�	QU7�$�M�v2ɱ�3��� ���؄5�0sűek>p=�;��2R�ѭ@���R�J�MY~�����95�m��rj�^��mY/��yOH��Ԥ`($L�v���3"!�5���#	zR�Ek����Y΍��G�pqs߇^�"^�OUz����a��u~幔՞H��ñl��&Rաu�#h :�Lc�򬙥rU/T
/��m�����.���Y.r`��"4o�h:+�am/c�t�׳y
��ﵧ�΋n�b'���������G\-��v���4M�Wz��?��؎���Ë�υ�:=�ic�oM��m�N��G#^p
+S�7�I�kx⓰�D��$U���}��2��^O/����>��~�'�$��b��y�swCH�B[�+U�(B�x)��ݨ
�W��<�LK$Lq8�v��/��%�����AN ��Tj%Z].���R�μjN�V>��kq"�^�q�+���Ko�[�T�*W����5�3��e��IL�,�͑
5�ܯǕ����D��>��\�ؚC(V�[���p�L���m�>N��T#o�o'�U��`���)_mA��pKZ�w����M����hr���Ҍl��Ư&qx�`߇qo��k�I�������fP�k�|��%�����E� 鹽�W�IW�M��0��W�agJ�nwi֊b�!E;���x�"�O_g���L3�
��e�v�zX;�6��W�Q%gpQ�]����˫�#l'|!E��^H��R]i@V��E�G���,�"��%9���E�?��! ��;P-ϔ�����Npp�]YF<��PY��b<�vtO���^���[�Z��SY�R7�U���@�m��lFp��玬r ��/��cD:#�,�A��7�*h�Nm�5i�#�e �q[���N��m��-MP���$'f�s��8�<�7֦�.g.1t�T9�b����F,�������q@�Ȏ� �����iݎ(wR[�9�t���(1eѸ��[�S��y$9��f(��?Y������}i��s�E�.ԓ�����*v��ş�?�Oe�Mw�^�z�ۂ�A<���j'y�ڞI~���:4�g�S>��Y��I+��h��Hwq<�W��� 쇅)�2=���W�n`m�JҔ�x#( G8M-��Ͷ�̃E%ô��6�k�X���łe��LMiBB���5�Y�u�9�޴�r�M�1�A�@��qr�)^�i���sa�ACc�|.�O%*��d_w!�U:v&�)c�Őװ.t�;�M
�����<*ڬ`~��R�[U]_kT���}�ቄ��9�/�Z��=��(n��G��*���y�Z&:%}@Na?=�h�����a�a�"O�2&��%e)w�>�0̆V�õG�[T�b�^OI�B��;f�N��
���a�{��Ѭ�u�'h���R���Q�]�B���Еv>�?g�xW�b�/�?��P.
��ŚJ z�Iܗ��8gl798v�p��{~U<����a����38��$c� x'ߙ�8�P�b��(��eq����0{�������;�sn�[-���g��b���}�c�c�Ao���O����Q�t3n(A���z����z#����p$�����LW���.�ϥf��'���\���c�5���_���F�r�I�u��:µZʝk4L("�w:j���O��H-+bՏ�>=�S��J�k��J� NI�Q�VU˷��~�Zf�>�����_b���cs9��B�9��eہ�"K�C�`��?����s��$d�\c��k�`*��:M%x�㝦ܒ;n,���R0Zz��l�����J	�����R5��'�ǐ�M�{��
cѤN�>�_�Ǳs:�v<Y��7��ql��ж����R�x"L�3��q�>s�&���!GcIր�h�*���'Ez鱬z�k�c ��5'�|���B�fcA(G&i�z�tu�|�"cE4��vN%嵻T�3�����*;+����=��'j��a1R%ݥ��cMpt�lԶ�=Uv���MIb!�'u��<l�f[˘?����������'�<O~/$�:�9�ܤ?GDo��G�cvPw#�&Q;Y���k�Ѯ馵{��-ۿ�"��ڑi�����-a"�����xg�,>��ZڑSqt���p��<�͵G9� ���Qz�R�_������Z����j��?�5D~/f�U>S��ܝ{<�:<�h�H��b*T�1�ͣ ��j�,쯌�M�f�Ŏ5��{�<=�}��o�V?�	�=l�7�����r��ɱ��� �q��+AA��:,�2.F吕�d���'\Sߡ��Vn��-ǈNl�������]��霖FDJ��	0�r�"�Bw�������E��o��p���R����iէ~j]E��:�W疄!�&����U&`�:\\5+�=� ��x�,�d8��_��f�m��t�͕�y�I�b�V�Q�Y)OB ����r�N�Y����:���=1�)���gɨ�yBF��� 4�/݀bTR��qI�p�$�,M�A6�<��[����Y.����T\��-J��"-��:;��]]�\��J>��.�e�~H�qrZ*֫�:�]����{ כ�ngI���y�S�����H�g]E����W�ȨvZ����Yw�a�Z�*�����N�3F$礧r}5V-��c�U�dRz5Y[��� 4����105u�r�KZ4�h�:��J�(Qu��I6����������ʰ��خc�o2,E�w�M�f�tX�=�����p�V�1!#p�+!���j��~��@S@!W�a��?����8��P�[D�a6�SS�V	�/v˂��T��7�E��3���2�4�n 1�H��U�W�V�DD�BAɕ{�)�VQz��J��+a�2��JY�89��yAjF�@�&��`^j:CL��8Ѭ1�,r���^�_ژ��\���V� ���:�ʐ<�V vO�WDI����3�����z:��SK8�on3��ɧ.��ۥ�E�g�j�yt@�!����oA��ޜlȵ�Q���A��p+ylܯ����Z�^�L����M%��D�����k��z������qVf^��l�zj�H��9L�X�����o7.x�nb�2�_����r�~��nd�uu���g�k��<#�a7n��$���qm&{�c�9?�}h��VNH��>_��(�t?SQ��?�z�ʠ�[�?l�М�l�?����okﲚ��6�G����5��:�jE���*e0ni�����X�T��"D���JY����#2X!��T{Y���~�`� �|��Ц��}e�xo^=����#0`-�j�l�~����^�#��e[��`KG䂽�<N|��C��|�����/���p�f��js�wGF������#vC{������y��]��f��ڡuW4�M1��M�>e�U;����23�dj�c����%c�,]��}x�8�R	&S5��.��*&{�*^�i#�C .f�V~͉2�{��+�p�<�9ɥp������Pe��LEV������a�z��)��q2$���2���.��;�(iw~�S����q���׺f\�<�w���5B�P$dg�R��+��Paړ���G��$�p��A��e]X����Zi��1g�t�Mh[W���a�����*��d�)͆rܡ�K.ܛ�V�Ď���������	vb�3�������4[k�8�O�ٱS�a>C�f����}��8E��.���)Ͳ�&��:.c�O��3���l۾�L�6p�?ˡa�Br.y���L^|�G�۶r�A����f.�	>+�0OMHBR��ܬ����@ �Ɩf
`�h^�]5�&5K�{�����/@�В�=�_��!��������ɬ�.�~jHV�D�s�^3@�C�� B����k9"�@����2ɩ�����вFA`��e�,��d��zZ'��ڟ�u 
N����YI����ȯSC���Ѣ_���<�;M�g�Blh6Ƞs�MC}ǡni'�"�g|$�jO��hT��?!k2��RE��H��U�n�	N�nN�Ƨ��-����(	E���������%��e��Y���M,*+e�]i:^brC�B��5޽�1k��������zdx�$��%�6�fu�[�I��h�&��Yw�:h����R�q�X�
ŉvh.9MDb+���o������a�!�$��ڵ2��cf�������f 6�s���aMق��w�2�d������k�Os����`.�m����������!�2t����%nS�{9��J��7�U¾`��Ġ<�l��O$˼3c6����p�G�FM��TUTE?�vM��~���(�-��hǳȱ�o�Ƴ |�9����b]�~$���������1�$��>�����yL��7�_j$�;^EQ���)+����� &�xԙ�{W^��� �}��!�fQ����S�)�F�u8't��� !2+��}xK��ѷ��5�1y�oz�2%����*?lkO�]�m�yK"�Qgf��_����W����Rt���XD6fu�	t��#�)1����2$]X[���u�}{��3�:�j���П�W>�e�k�I�F0�����x���w��LR�l$?���۠���K���_�"���`�P�"����g����c�
�ZmQ/&ԮQ�P"��&7]�/�=���\��r196	�-����e��5�a�!da�s�|���5�w^���k �ì ���-=�䙊[��N5��un��H��1�>Ui�&q0S��4ȂB�{���w�^"�di��.��j�����H-�x�!�I�U�X�x����w%�.:��/�#^Ob�6<�]񬄨
��XJ�g�By�������m�+۬�wq���;��h��^R��]��#�����Q��+$Ů�)(��%�S^6�0D���e�!�]j奮��$���/�O�� ����rS���(���t.��o��@_���4���Ue��h��&x�A�n0��������]�,6܎m��w���Er��&�R�\�RR#D����oh9�D��W��M�>3��U��k�F+X�^Y���-&=w�y#�<�����:aF�g�j���|	A���`ul�����Q��t� ��)��l]�̨C&V`�6w�
���f���oz~(�^L�0��\x��ވ���,vt =�8'�>`]�wp�VU|���eQw���m�|���z,( gd+�}j}��!c�[�.��w��s�2/�:�~��&A4�k����tu��0>�G�*D�՞��m.�2s���?ӭ���u0�Y'}��yɜ�h%�i�Hx/���=�)�OV�D���I���k8�P���>�a���S�m,����8X�z�����\�]Z�=����u/�o�ȣ��� �y�.��&��v��VBt���_;���#����F��t	�y�Yj���M�zM�5u}Z("V5���s���զG�^�:3��(�M�A���P�$y��o��qU�Q���y��d������j��㰷�د$��/z�<\��.��p������\��^� �"G�A�2�����B�u\�D�U�}̓�L=���?��|��-��[`	͍��[���r�~�n0����ߪ<o>q1"\�v�j�*[�����E�y��p�1�$9�'ƩN� f{y谺�X#�������y�·��7��-gT�c1�Bqg�;��hc��.��/�<8KA����둦C�@?k�� ��G�o[>8��x���F��#_x^����,t(ǥ�˛�xƅ�?��`�r�h��a���d�>�h^̄߼ȎɅ�p�8;�y� ���b9i{��
.粛����U|ykڢ��$���[X𥄊!KP'���_E f�֥�?����t���L'U��:WRh�1��]l�6��^�ʣ�U��p���nG�x�S����I�͎���j�eE-,7�D+9���n�
��zd�ڍHK�+�j�f�*����A
ѣ`g����H��ZH�u��g�aؖ��j?��'쫩9��j��mʛ�Y�����f"��~Z����֑���9��w̍�BH�ʽ�3�Y���D;���8,x�Qj��sZ��+o'#�Lg&�V�@�$P�|��`�ߡFRaI��㮜6�j�N�B�p2k����;�I���t�5�=��<�e>RH�P�r��W������#]�J�4R[������i�I�o?G�ec�����2i��?��s���K`���7�"Q����r�}D+X��=6�޺>�
U;$hR:�S�٣�*O���]�AB�s���)�:6�����tx<i�\�VcѸ�I�7I���GE�dx-<�V�@��1�ΪO�ص�����%]�c�� }s�/���k�7�9|sN� ��<���S�ǵ�Y_��
ݦ��5�,��.�wag��^�����?}��hoi����?�W+9�nU:UM�3ֿ�֑r�Rb<���X�����4�
�)����ك����A:��x�������S^ޱ��؍�z�vc-��:[U)���G��^���C6�Ү��XC8�R�]�S���d�@d5������H�
��*���Z�ҥ^t��| �ޘ@I%:�^��Eo��7'l�co��<4�}�}GY	^c�1*���P �6Gʋ����h�G;,̱�*/2���ˮ��L���-vp4%�#��9 ��(�a�f�:��ڞ���vL������I�Go�f��M(;�FNt4}�a�#��Bg�5i��,��~}R��FF��q&4Εd>ۿ}�K�I���ʙ��./b���b����^;����}��;&�tj��|B��~�)[��[4J�1�ۣg)�}�<�4K�S�c[8a���q�3�8u	��Ӗ�wc�$��sB��^�5�����1QL����(� A��>�0!�&z�>�����d
�9	�i���\�U�.�u��W�>��Ak�l 6wN�Q�-|��n<l��SS�7��������.�܀�������g ����﹛���hR�R�]� �M��լdD/����01y��[=���@IgCy&ޕ6���	��lv�X��*.k�O�ŪuJ�l�hb`��B2�)"�����cxB~�M�;ȟ�rx�G�7�<��,V���*	�dH��4*�|�+�G�%�"�w��-#3dۛ��ۑ?JD��~�+g����L���v�D#����{Y�� �{���s�U��?0=��S]c�h$0��H'S)�����V8菓�q���Օ�m�m�����PҮ�&w�����L��I��U��$y���^�0H����&� 2A��)sb,���Sd�n�C/��9}5:1�r��ƥ�|�,n��*��r8���P?�٨����M���p�DE�'U�$�|����m<�{ȶ0P��-�f��0ʟ��~�D��R&�P{�Ԕ�{��]\9Tj͹$~ �Tw�:H)�1F>w-�3�4��/�.�n����. �/B���1 �l�m?*�J.�8����{�1�f��3`ֿ'���sĔ�ŨV��g]Q��~!ӖH�j�Y��.&�-�7	r�q��~���.���k�(9Z�>=���(�L������+�fh�NI��S��7�	����/����jh��2᧿�H"�6~'�W�����b�%pp���i~�a66؆"Dq����%�`�z,i�β8>kx��4e�#Q1�լ�a�/���F��d��z\e�
��a�K�5r��K�,�~�E���X���u[�F\w��Iﬠh-B����͟h��v�xjY�_}����%���0( J_b�TF%�+�l�q�
B�	Kt�����S0�|R�W+��Y��O��ơ��<.(S�u�A�gi�&o�A݊e�Y��� �n�pB��&َ�����;v��.R�:c���]����Hmm����������ڨ��ҧ����ٛ
Su��>]�nc�&8� �s��F���z�N��V�x���Qfz�����@U���6е�Q}���X��
�ٓ-���:ƚ�*�p�ɶ2s�������:#H�- I����$�t��x�@���T���f���am|�u�uɭ���d�
쓓��]��.@�qP��n}e�
�d<D�&<��=cP�+�P��#j�� �S��ޥ8�7���|�+j�6Nj�����R��q�����1+G�w#����
;�.���rn{c��Ƹy`�d�DI�z��[�t�9�K]���J6J`��O�P�q�]&ng��/	-��!kܕ7�f��S��Pk��SR��W�U�ͼ8�]�<�~D%t�L8�P�7[t����[��|l�� �B�#r͎�1-tZ��8�lP&��{�}���߉�'��X<Mm�]K?�a6	i=��U��,�3Pl�)v6j5&��$>WϩT<W�,.b��'�x�"\��	K�)�8�s*�H,���g9�p�7���@�H@�RtKᦍا��`��u[��]�[Ʃa�spf<̴�J�s\F:�4x��V,"�<6{����q��*�WW}�)�����}^���J,�o;c������!̫�V�@Ez�pAi�����oΆ%�ȥmیg&è)�1�5Y�'<ő�ʑi�����A���8�+gw, �?�㝠�:S�[D�v��`\��DJ���r���ma�"��x>�t��L�ފ���Ūy��������&��xa�Hl��t��y�50��,Cү�Kb�||IT�7�!�f�� xP��d�\�;6��pŒ.wݒf��[���"x.�;n��~pE<�������/ϓ��)���4�����nq�,���������,����oK	� �=l�Ci�L�Nٍn�z�r�ݬ��4y��p�!v󍡵�=�"�'k�8��@���~t���[	�C�Q��^�ct���O�U��>���$	��C��#����mG҉3r9��Aѓӈ|�i^g5̬v�[>����__�pw����V�UC�k"�]³�a��7�`�!!k�4\W*���vb_�}=���\�Oa��׎��n�z[+�w��.���y�-��LZ�/#��4^b��?��ƀˠް3Dg�H7���h�;��z��Ж4NmHRVC� ���v<���� ͎��l��o�K삵���MC�`8z3xW��ֹy���V?�Ea�R�אD����}��N�W��=[dW��&�3�Z(��7�4�!yW�e�Cl�f\�WSb҈���Q��9hݓ�ީ�)Y+��-��P�ς=���}c�`N9�~cb�]�jE��AN�j��1D�O�|�f__�������{�{�?���KK6�
�����wx �"z/+�W|�ڒQ��^�~tlC�(�xq_Ke�1j�:ٖ�ޒ��'�f�XA|���)$�4�~����E�
߇��&��%Iې���v\S�RQbnb4���y��6^�g�/����!8�Q�1�"�]�m�.
{7�����j��Hrz ��B��O�i��e�4��s�˸�e��3�z�?Y'��C��E�"q��- ��l���a����lb<�U�)4vФg&B����א*ԀXuY��>��;,�fe�zW��b�1�^��WM����>f�:�C4��?�h��!��}c%��h��:#��F�V����g����p
���Q2���b�D��f��$��#fpm ���H^n����<ăs��㈷�6|�c�R����P�?�Ê|�%OD�2lp�����¡vȮO�j��q��m��u o���<��SCVԂSy�,s���[ z��S4\��s��~H�m���	5<�ɴ�O�7�9&�%)g���O�B�ઙ2)�m�pG�3Z��)�y���3����Ꚍ�@�TG�V)�m��̞��w�z�W�p��l� �UZ��В}B�Ɠ�%#:�:?��1H���΄}��QD�+��!�ߥ��]'��w��V��_t���N�EF�C	�'��d&�y��J?��F��nS�1�RR�Mk��fA5ɀ��h��x �����i�T�?�!1
G������h|O������C	e
�Nt�9�6.�� UD0=��k�`A�*�h��"�Vr�&��4 5�6D'��+X����"��g|�����L�j�$G�ݩ����̋G�V�b;�=�f&�B�([ep�2�P�"�^'��C�qSQG0�!��?ks�����0wSI���������+����x��[ܫ�B����(X�S�{M������/R�Mc���Xm*�7� V��9���&��Z�wЙa?&��ݡ=� 0�ĝ")��xM�F��QQ�qib'[��"�;/��P��\;�CwB�k2��1���X�Kʠo���q�~��%�D2�M���!aĸ���?����������^|��wK0�C3HO终�o��z�(�b+R�Y��f=ho�#M����ڟ�i(o�j�3�A�́�ˡSw��xv�4;w���{���3V0P�DG�w�#�|%�F���
�6��ot!f��lR�$K�ڈ1�?a��rb�J�Z�����P�Y�	����SY.�-�!i����%k���~ja�E���x�a��p��&�n���\���&���z:��5���U�E���V��V�T�5�M����V���Ꞁk�qM��u��l�`����uML�R�ڝ��V�lZ�*����n��5xb:��f�@�o�B�)OMQ�i	B�,���I���1 T�U�C����mۆ�։XMB=0|��F�f���jUZ�wNz��&������LHN:� ��!�OH
ؔ�,�p��`��~�������xl��;{��&1BC�H��_��V��ӽ�|Ԭ��|��HR��B�vS!,�u�$^wlGqU��ǻ�x���rK�C�G���F�<��(X���H�P�RL����>�k�w���s3���d�I�`�.)RR���A������x�&B��e������C*U͌j+����A�\���G�����[c
[l^5���ab,��*L���=���lynj��^��C��r��яv�z9!UWN���ܚLm���L~i��N���i����O��L����	Jǆ~l:�^�6.����yD-�(j ���Znk����P�[VB���-�:y2����&�����E��o���w2�c%E겶��q�z�|�e�~D�f� *�����$+�TZ�:���3��E�{hع����Q�L��[��Ԗ|<G<dFJ��Z� ��l�k��3��Qf�C ���Lof��-��C�����ZH_�Ggr�%!�d7p�6ְ�g-�]����!�$\�Xbg9�׆U,Mv�Q �j�}i��f�A��g!��P���	�=���^����-�	��ɡJk<=������m�\|�og��g����!9��%+�'�VC�Og5�/��d�l�y!N�RU ]7`�)+Lq�|���>p�<��zI�.GJ���ۀ�n
�V"��'GS'$2���H��i�	�m
u�]}j����ّ��)V��eA2`���X���k�r(�N���M�O�_�r��S�JЕF��8YL�Ȥ��k��ak����a}�*qPKP�^8����v���Ò/iU-�-w��"f��sĺ���­Y��!�u;�"|�~^�>Y���\V�?0�p�" ���y�G9ݲHM�� �t����}�(�8�������Z7��ck2�H�Ϭ������[��|�/�m�Ҋ7�u��qOl S>џ������B�P��\�Y��|n�Vu�ʽ�:4�x)D�G����+^e�����ܛZ���Q���_�x�,wK�jN��n�1��o�P^abs�{��������a��<��68�;#�SF��'�ó�oBF'!RcՌV��)�5ᰧ�5vQ�G�.�Xz&8�zחö�=�bgh:�-�ns�1Ƴ�=����a[d5Wyn����k�ӫ?*�h��1}SF���Kvl��M�Mٯ[�A}"]^	��>N�a!�{��u�o�Je|�he�:X!�T� � �^��c��ė�Sr�S��Бc�_K�񪡻�On�H�K����3`�c� �i|I1/�@��[��Dƚ�ǿ�����W�R��n"\]�m�f�P��?�����?M����"����pk�\03�,�� � [�����J�)w���d|`���Z�2�y�YT�4�",
�;]ҥMDyL��k���0��q����ه7�!L�>zu̱�rV`[�i�,S�IW��80v���XR�9��W\SHFIT��Y2�
�I�1�J�V�NW�Kd?��)����n���
7l��.�^� ��6�j��� 
�H+:?�����X���(�eN���+��ր����KE�/�X~�X7��b*�P��u�cy�A{`g�1�"Ә͔Qr���EDC�U�U5O3��mm��n�/<j3�{�Ɲ�C��K���U~xi\I�����<��+�GDk���!a\�₈�09�r�I��p_�+��HP�o��5jF��PK8ܼ��R7�}5`����S�xd}��Z��END^(/�Dh�L���Ay̼�5�7ɋ�"��-�#s2}�K���`��Rv�+��M��W��m���6�;�5��Y
��P#�+B�G:��l`)؊��1�	
(4�_F'D�G��B勶8���� �D��t=x��c�1TQ��[�q��|�j�Q�]�Z���T8��cۦ��By�Y�>m�S�Q�U	�Yl����[�V��ǳ�raf6I_O~i�\`9-L��� Vl�H�'v��ЂN�m����>�����F�"�<G@��V��:��a�����0�����.�;2�]�A�[T(�?��2׽1/:��R�-�ޫ�1 B�;�y�� ���`�cf���9�K06�-��A}�lS_V%P��ĞB��K����D�^�;�(A�	}2W6_5��<7|�uqC�_K.��5����B�ب:>��^�}R���?Y���^K#����E���޲a���;5�R����z
�^���kh�f���������Q��)���0�F���*���d���:�׼���0g�������G��̎�u��%hU��g����be%Wve	%���va���p2KC��������tgs�4�ws���Sw����]xx��_���R�����]|���sUZ�(7�rj9�p� \�>�oo�d�|��M���'t1��OP�E���}`�SG���%��dG�	ت�0e6��V� \����0��r0Yb1P���1�����+S��-E�`�,h�2���&S�1���I}p��n�m����o��{0�#I��2���eah&X���!�Q �d;�{�(b m��#�Г���W���	
W;"��2�P�#�
0�_�:���N,By-�;�wƇ��v�Ri�CqTc$JA��[q�v�Қ8aЏg�W�F��[e�M��C<)�9��"`a��Z�E�<�\{:?�}��K�H�;V�U�Wyh���5K�ou�B*0f\�t)�<�<}�
����-W�L���&A���Vv�%�����l��9�y�?2<����pd6I�O�h��0����N}ˢ:�� L,�#����?�8$ML��*�v�^SU�t����p$���e��F��,�Z)��U���T���@Sv���]  +��,�f�� 8���yO�hIOˤ �B_֗8rH��E�����X�K�)����Lׂ�5ß�P�t�,Vr��:�,\�*�C3(���&�䎲��L~�?�}a3x�Rv֥�|ʪ���T�ltCcUz��h'
�eOR�x}0�t��'�
|m�%X���%�tE����9�C�Q�Z'�b"W됤���5c|5�U���xO5ﻸ^l�),��즲��~
��zZ`Y͈]ϊ��*�k�^��-��qY:h����d˯��]���M������Zܙ.��!��N��=��e����^���%|@��Cħa1`ث��5�Q�oq����ƿ�g� ��΋��E��AreW�+�
|('�*�|�ٖ��h�;�������>��˯ ��B.���,��iTk���>I�Z����l¹C�⹿)�M�|���۵U����\G�}�=���8f'���#}����qIʺ|Ī����l[����k�S���}�f�P�m�C��i)��%'ؾL.hlI>�wF���>���Q*y��#����Q���n�+���H@Eۑ�FC�~}���� ����U�M
��_��.+��&�B6�y!��$n�$kgE�x��]K{��)���L&�%N����PV�����h�^,y�܀�/��7��7����=p��	�q�"W��}������<Q;\�XH��2V��Q%�	�5���JA����t�E�������ɠ		�/�~V�zkL�5c�X���5�W�Q]ͬ��Fy,�������~�>�iR�� ��I�NL���l�q�g��Jm`X�Jک�x[c�r�Dk ��K�*cRM��`E��=K��Φ��M�������c�Աj���-'������5����=Dq���r�b����ab^��$�h��`��߇MmZ�:�B�����	�OpC)�̟�o�6v�aǰ�e�Q3Z2q��c��8���@��h'˓�zЛb��_5)���G9�����'��r1H js�P�撃 �!�j*�{5/K�UA}�L��B��Y��p�\eĻ�B{�[6�e���As�&�כ���qv�����8.�*N/�A��H���u*�@9^�\ft����Ha��m���E�D����.�9�Xm,-Yp�$��g%���W\͖I�!�VAp�3�W8��ٯl�3G3R����(� 徦޵ȕ��phL[��?^�?�Tf��+�Iꏮ���4������i�P=x"�Z���K�"R*�C��W����Ϥ������l�V~B��	�$�v�њ"�&�w�Q��0,�vJ_g��"��II��O�ie"��7x�1�~R�@��#�����,��"?yV+�t,7+��[�	�R�nЄd��O��Z���p+�e��>�m�	]̡u� ��M�ځ6��É�&���O�õ+��gqR�Mi��E�?(yO���miן4l����Acz�2�r\��_���ac �Bw��Ri>��K�ի�C�%���u7���,���S��k)Lf�6c0��n)��\sm� t`�Xī�Fj�j����7J=�cs�����I��������!�T�X�K���|������"�_��\��|J�v�g��❤?�&䫸��9�F�7�0?z�[�ΝN��P)ɛ�l�<�t�s��VR"W�0E���M=䌏ˇ6L!I����ȏ�#;Y�2g�z*�������\H.���bh�E�%ԩ��W��h�Hjĩ��a��T���x�ƌ�/� O���]�5�������@,�>9���yѹ�n��1�@�%��ٸ�+�M~�c�X�J?_���;�B�[밳�CI�(�6�s^cvE `���pV)���S��:ֈ^aG�%
�����o@�Qij�g���Ʋ�g;]��4~��J:+;T�ʼO�˯sn�S%��iL�@�]<�Bu+`/�}�h�ّꁽ��\���<d2�_F��w���K��ж���|+M�whO�#���������Yh�n�3� 0�	��JC�:0�^As���T�\�'��:��BI+[UE�MtO������:�ئ�b�E+'ê���s�Og�_ǧ@毮���2���w��ʔ{@��w�y}�wIŠ�a��H�t�����l�4�0d������`��~����>'p��� =�P��]�y�����	q/�.�O.�\0E�^���ܮ{Y_�Xi�i:w�<BZ{/�
�|&{�#"�F���l��aq'B8/�����ZO#�s�u�4G�l``�@4�6	�����J����86��Ff�����I��a�J�ғ��0<pFů����Q}r+�9�)�f�e�$���X�憞�ȯ��/���v��&�C��8H\V�V����L�]Wu��t�a]"`��.�;|�V�^���c�V�2*�ٴ�P�N���
G����c��զ��0�?��r�V!YP&6AЄF[�QJ_�e|�.0ADM��9�-V�o�Ă��<G��_��ō�o�8��Vl�ի�KRw�ޙ�&���4��r͖U�[A�Y�!��g��!j�K�W�
�39ٓ�D�qs����4.Ѳ��|�%дZ��(��T�t�7s������^BQ�c�	�Y�u����a{��_a��\�	�A���m�-%�0%@�άnz�g�iF��V���w��ۚ
߀��R�cSH��#�SD`6�4� PR*�^�T��w���;-���*s�U�`!�Oa�p֮eh`�a�z�]�6����эAX�t���pDt`f�����81��x�Qv�۸)��#>6렯g�b+��'���?q�VZ#\[ ��>l����J#�m�H�$�oq����q��Q/�I��8�����z�23�(�U�x�+pŷ�L6�d̐M�4z���X�#_gՎx�c���;E"������?}Ոn�|2�<V\��{�3/�E���ф�P�x�X�Z�Ň��x�=p�}{@�E��2�Zd羍�5�g&Rg�����K��b�U���۾���^f؁U8�;�B>�nwI"VћS��7խC��l��z�����4�H�D�I0�]�eȰe������(e�sa���B�dj�����M���>C�O)s9�n*����׹S��L��3��d��}�_�O�rTn:��<�jn�'"�i�|*é�w��3xj��}�HX�T�2��'
���s#+�y�O�+c�D
䞮�s#H.V5.�L�Ee�돼T�(3ʳf%5�YRe���Rk�7��Wq*#�M�.7�G�ᎋ�c��S�n��1u����~Ҥt�(��y���?�ء�Y��$S7i�� �^	�Q�CD2�� "[�1.޺v��k�"�佑�R�Qj� ����/b)��Ѕ���Z�;Hcn���<^V�
LJT���t�}Ӡ(��%���a*Yܝ��H��������zy+ �Ĥ>3����5~�{0Wf#�X�Ρ�ԥ��ԇ
���݅��.���]w�ڠ`�22��:���I��yh��k��Go�μ���O�tng�Ο�#a��;t�D��N�h�Ç5@�4��mÂ⧶Ǡ=�2צ�e�^���N2����F������4��3���\6���@`���!㎿c���lԂP�������߅�ȴak�5���?��.5�a	���� ���Sng��-�"ޠ��g0���Ж�g�z��?؋�c ���d(���wd$ �����z�k��5��[�W"Du��P�1V,�Ze���a�P*����.F+�v��̤`b��c�e9�U���{��L��B�#�r���>-I^�d۹3[��ǟ*Y��TL�opw�5�x&>�̰5�)dd<�Ar�����u~��z��wg��µ�4��pg���(���sm|�w�mT�^ ����$"J3���e����B<ʅ�>����"�ڙ��D&O�R������:�h˞)�MAc��c���	,�:�9P�?u�W/�ӾwŰ�G�{'�`�s�]XE�{��3*���*���**:��q���|!Pa����䫐�	���u��,�~o@�d53 �no�<z[�,���M����y$�/��P/d/jΈ�y��=�y�U�ho���y��>��61P'�WF��E	`9�n��lg�����|��mV�Q3�+��E �J;��i��g�oϊ}4���[W�r�ga�$�01��$d��!����%<�&Y
%h~�߻Tv���bR)"�~c���B�Z>%pH֡�P(Bi��f�#������kSx�m�Ws��5m���Mvν0�4�*�sO�}��o)��m�$��#�J��Bn�&�z��ϔ�[0 <h~�w�^Ձ?y��YT�(��1��7핑��~�<�Y�k�+^c��as1���Uv�N�˹��r&1E7��Bv���5��ⳟI�TdrS-p��`�����^���q��M�����P�'>�N3�E��m�(Q��m�"��V����ٙ�D~G�+Xz	(Z�VW�JF���#��������C?>F���R�m�9�6 1�A�U��כ0���]O�
���vn�:D;�����e8�V;��2��4�%8çV�����+�9 �5�p�e�<vO4��G���=^�49�ݠ�	0Sϙb�T���)=������/�q�H�%a�r��:�,B��B�k�!mŝ4�id��J�6�	7�)���������Z��O����Aj���'a^�(��1
皭{�,��7c��n�{Z3j6-�-�+�����rR�|��j�jZLC`'��]VG������NL	���\tY7J�q���D �,���]f���0�N	xd̖V#OV�ϟ�}�=�wN���D%���?�qa�oF����C�l
=x}�g%�f����=0����5����C�{��c_����7oj�y:�:E��hg�H�/jqx^�"�	3h�LL+6%�Tja�i{�5��v{�e��y��>?="�s���b1&N��A����UWf�@�H�}8U��h�l9\�૫��D���?C���2�Q���=v�����l<疷{{�0x5=���̷����ҖI��z��֙��Uu��8
��.i���"�_l�Z�!1��݋�eƬ,�l)���������M�2Lvh����E�zB���J�>.� ��Ԭ2%H�L�$�y֞D�T6��Pl�ٮُ,f��⃱UR�������J��W�я99�]M�S���E���
�G8�p�/?��Q0�k�s�D{2�$�:g����L�Y��}�=TWV�-�_�UC]�>�ꆱN]]��K�-��l��.|�#�gMy6�s2�8Ĕ��4d�@��=Q�}C��i
6JI߶�)�sL��� P2��h���Fr�}�e�h���dc@��nyL(Su�w�d��}��R�;�Ӫ`F���Ņ����o�/���f�����6T)�,x[Ia9$8%��c�b��=�u��dasT��Ð�8����Xn��n�&v���g5k/��;��gEt"T�E[52�@[��^j�Jb$v��q���������9�q�u��(�YvI�T��u�*x�pS�҆�q��ޓ�ſrE�W��@�+J��,��QS��2�!OoϚ��_�?��>�E3�V��앆Z�'=�\��a�K���������YA0&k�.��Q�4܀� ����WK}�Q�p�)X(0R��n�z�G���]����ߴґxSj�������Åw`q*�MR:/�����a�f�)��?.9�	�^q�&p���f��2$��Ÿ�?���O(�Ru��A�𢄘���H�m+
���#�������:ׇqb���9¡��\�o�	ѧ�}?%i+1�Ia��r�$��+e8YBK��vc(����s4^j7�?�?(2�ŀ޷H �|w�s�vjwP� +�8�S
�v93:%>��:�ƀ�H�ஸi��3�M���A�ɩ�ԣ���Q�Aǜ�sb������p��fcri �-Q3�;���r�ӄ�����J:��2���Q3·ݍڍ�1�!�A��+�J�g&��}Q�X0�鉳�H�f#���y�k�����zyez��U�uN6�rv2MM��"x�M��x�X*d ��d{q?LU1F)�c�\�zalw�����{��C+��Cڡ>�L�T�d�o���M.Y��Q�zCq���!a�F�#]�}����@������3�r�}�V��u����TM�M&JqxJ{����m��Gn�<Qʧt�2@n�.� !\�!�(KW��뺇&=�+�*)۬���S/���A���~�Q,z����-��WE�S�j^K{M,ޏ��A��p���$�����ߙQ�C�)S1d	�4���(���M�İlG5�1MY���H��(�p�C� ���ת�����ճ�6(�}���]�TŅ���5YO��d��S&q.��8�[�hgx�>�9���8s�ZI����ټ���҄U �X�K��Ew%��l���f�\.�zo���׵�d�8���-�E�J�6��G>�ȥВ�l7J�?������x1�� !�YLI )���ŻP���YA8�"�Vh�V����~9l�@pi��3�Ɪ�C�KI���JYW[�vu�+s�h�y$��T�R1'�'�U7ry]�˿64`��രN٧m���7�:1�E���ك�ŗ}�'����(����jbuZ�]���ں"ȬX��m��ˊM���
�����S�P3��������X�7�k�%F}���������B<�)ꮗR� q"�K��smN�>�6�F�?������V����a��g���d���d��ߤ��Iӿ��f��mZ:�L�<�[�=g�=�������3� 
'�O@aq��;A�W�?��<yn�*���7l���W����e
��n��y�_]���gݎ�>(W����x�b��#*#�6H��1�V=�Ɩm&�c�O]� �1�*�#Z�&i�8S���:=�� �71��R��,�l���2G��f>�B����6�H/EA�G�]A�0_���X�6H$�CU��S	2�|Η��~�d�q��x��V-��$�J^k�����%g�G�s?W��:�ɴ]��a������wc�� ־9v��=h��'V)R�� �-|/m@�j<Zf�P��0s���:��!+�Ԍ000Hh/%���.P�5&`�۟F���
���魸!�b�*�E�P�,m����J]k��:���"��55A(�d�+vvl�_:'1���R����uR#Z��2�_��(�f����~Q,��b@D�^n�X%�H&2��s�͂BiQ�6��7}&��z	YR$� �l.K�e4Ut6��l��M��ꍓf��l������C�`��N���JUv��z����x���������Ǆ��wg�
+L�+n5	a���+#��k߄Y�Idz�KB!�1ɻ�eb"=����V���E�bk����u;�5�ћ�����k�����v�E��r�;?�6�!�<��X�黐�|I��|8t�o�c��׆�3�D��eaqg�:)1��l���S)C�b�e)�u�g
�Р.�j}��q�A�r��Y�͵q/���e�܊��F]+�����ǧ��Q��}�H�?)TD���-�!A���"$c �㟎Ϥ�!�@��OLwiݯ=z��4Gu[��#��f��e�������5��d�RCЌ-��'�ow�<$����c��l�� �wd�n��<���0��N�b$��-Mn  ̤�z!f�F�ZF�C�,'�"�R��Eε�1�>T�>��^e��d0��M_~�kl)C�������g� m�uB�b]��	v^|'��J�KT͂�Ν�L�t����(d�ϵ����v���_z�$}�?����4��î���%ϼ�y9e��t2 ����a}�Qx��\��2!Vd�SeR�q��DN�%
�������L��a*^,k�'t|�b�f��Bm�=��x�,*��R��;ҙ kb?)g�L򱎊H�@L�:��)BeUt,�N%� C+�^brE����y�ӅAAUN4�FL���uQy�㧌9���� a�Fm$`�[Î��n�9��R�����������։�Ĳ5c!,��9�D2ЧJ�f�9T�ŏ�t�\;bn�z�Lֳ��K�'$�m��/�>�C�Ж0��9W��i�W��F"E(d�ke(�ZR�bTh�tl,j�"'�T��
��C����W�%JKͺ4��E�S���c䓀aQ ���6�����zu���t:�$R'���iIW���]�^�����؉=IUwf*uƤ�x�\Tos���zV�jM��#��
�m�Ѝ�m-�L6�K�;���>��������sn����
�֊3 ?>���0j�6uC���g�ⷹ��1�6�>3&��\w���p㆐���k(��y�J��d +������I/_�׵���R2�ʞ�*H���'�x̹t"��C0n��K�3����/���>u�E�HPVyZ%�H$CK%���P���ei�\0���+i��{^.��v��x+H�k�d��ɛ�`�V���y����'���)PWl<��ݥ�,��mvǆP���櫳�U�y�}_x$�[S]�xWFKN�����y�,D
U���_�n��I!Q�Su��pB.�#�m����!,<Ϙ�[�tH��Vn�P�k��B�
(�2�6�q�k�,HB�� �*�CCsDEޙ�s�x������H�P��T���
��j�7�)���m�"5_c��}�-�ך 6C��;�R����E�F੽,�m��N�t���5����)asd`.�Aw�i�ugT9�g7C�m�m�Ϳ�h5����!z[x��!d"��f정L�d%�mrz���/j�$�B�y��B�ح|@��'�[������3��k��.!n�{KSPf;Jݍ��_�I_���D]�No��N�S����.��Mʄlz:B��/.�Yr����Bb���%z��\��4+�S6�R��P�t��HJ�ፚwiȈ�a�����3���V;�Σ�Vp5;pVl��������]�:߾lhjt�|�C�3�AXd@ϳY1r@}m�a*9ͭ�8����P��d:�D��lv�g���bqoL ��_֒TKw��vxA��:y;iF;+@72�Z�uR,T�N>�tb�
�L��ӟ�B���
I&$�z�S`cj�ac!��Y� ��@���ɍ$��؀�j���V��#N�6�\b�"y#��������^f��ǽ�<Q-&��㻅F&yYR'���.�F���+�MZ�P����O�Rr4��9�-��|�7	8��Q���s��J�Kq�m��g��j�l���5)l��`��E����k��A5[5���5S��>G���e ��
|�*�f��}R���:=���[�m�c��X��ӕ��z $1�~ʆ�h����U��{��3r�%�sgB�)�E�U�%o����Ł^�	��Q�8�˻�b�&%10om��J]��C��p�^�e6<Q��� �g��R�T���#�j�����T~ςq�����':xG���{D �z�����˪T���Tu�T�n+.��8zu�?�cMli��5�Rs�k�(+Ak3�|�VJ �7��ۍ��EJ��^��M���Pg���\$�%h�Db��̑{F�z:h��بߵ��f�'	�!��[kh�v$�>��#F��U�5͍�^`㭧�em��v���x2�'��UVI��r9E�:Ew
�"Jh����7Iw�$Qm�ǿw�GO�[����-%��f�7ق>�2��8�G�%���ę�#�	�5%��P�S�b�$�ar�������+���E7��0��R���.��I;�.�P��*Ts�iB�L�٥ƛ
�VP�{t,�������c���N8H����F[�Q��.�6u� �d0�P����rzL4s�gE�0���9%���=�9U�j��:�&>��_KC��i\��b2������2Q�ڌR��Ϥ��@�I(sڝ�5U�J'�?6��
�2`R�C�\���I7�m�}�Um��&޲_��is�_�$�2X��yF�F�d��ՇG�l�MG�h+�j��ix�I������8�Mu�q=�m��XeG&r���A�p��~*��Tۚ	 ��JD�?/�L��fH�ݘ-�7�-�5��td<�?�:�g��}��N=��;$�Y���K��a�bCO�t"{mE;��N(~�6E^���4�\!�@�\�w�����\�)ѐlQ��?>�~pu��y9(�>��r�?;Q)����Z&;wc/n���<X�|w����H��e2�O���u3L�pRc�k�Q�R9�p��3��x�{� �Md�Q�t� yv�0�hjH�U�e�L�f��#����@	��t��<�`��]�#��:t�B�a��R,�F���Þ@���v~/0K�u�Q���\�ޯ�^.����D�-���LGA[2@��^�z#�#١D�.�8%В{�[��GO�m�J(dj�����J'y�4�Z��R�"���It<�">�F'Ln!Ҽ��>%�'�R��nlv�tT�w'޵�I{#�}$!�,9�����%|(�R�꡺t�Eq?N�R�&9���Wk2�!�����(��a���=)Ê���?���K����4��_�WR��~tYʳ��R*����q��ap>@ �9̔����Dܐ���a�B���
I8�J��-d4�^w4s��H��M��@0�V�p��)"j�1|DvZ�I��>o�
U&Í�G`Eǥ,C���7��9#��D^�<�5�y������,��?y�WMH
8�r��}9�4=D?u�����2�`̕��PGK{�NU�l?*���5��Ja���H���J��Q�D������6u)�<fPsNB�9�AA`)D��$��#��$�t��P��=h�2t�	#�Z�4�����6/���ZXMɍq-����a�@I�a?��϶�s�	��B��"y��R|��S+JĲ�3*:�RAd�,y�����Lպf[ʔ�*��t�W���#�G(�w����'AUnْ1:�=0�Ƨ�����~�H��4 <��{��E���^�Lй@R���a"��q4ƂT�8CT"�3�u���8�k�@B��a���
�<AӓB�Ns�	�W�B}p���w���F�i<`�olTw��ݡ��Ӧ�p�O��r2Yy�)�����6=�1�4M+�zpj�UސH��s$U�S�z�:߶je���L$���t�� I&�wW��X�)JeV5���bG/4qv0�����*I��[I���rWb����ᆉKh��f,8�K�"��6(�W5+7;YI����G�1�2����]��L@�"/����E9���%tD�<gN.SC����C���	��-�ϻ�P�Odw�W�|w)�ĮK�+$��îpȇ���6"<E�j�S����V{�m^�34�$���s���fӬ���;�V�������b3�vw"��q�"~쩉���<t���|��w��-o7L
�մg�!��iO�tk%&�D���܃����l�b��2���q����)S�Up�Sn`�5��	���1+B��������,�gK]�]��	��)SN���]�o�` ��b���?��v�f���-���c���
t�Fq��Qد(�,%	=�L�r�4�Ɛ���B��13YU�`c�D�թ��-y��#uK�&>z���"��5�ٸV+U���(�iAnJQ\�^E�$�b���(����OO�(Ѡ��?yy<ŗ(*A��䢬cz�~Ai���+w�ռV�(�A�7�2��f����͈c9��ß������g�SA<��5V3��Z�Г�)Ű�X�F����i]��q�l���I���fR`!8܅πذ�[��,�¯vġ����r���qeƗg���˗*M���s��Rt���@�@�ࠖ?��x+���\-{?������Ή��Q�?�#�4�}/���x��3{�w�-�!�� `����m��W��y��$�����R{w���_��ȹ�H���[A&�jk%>+��vɕ�V�V+��.P~��\	Jt����H������y���d���a�F<�i+<b:e����>�mE�U�r3��9(Z�Wb_��I�Ky�A>�0e#Dߤ�b�^л?���c��eae��7_����j"[oc��� �9/��WD.+���cR2����MtI�ؕ��z�-�1�
�t���a��i�h�k�A�nU�bl�d�������b�����{&�b�Z�t��������u�M�vC�����J�i]S�)�"��z�䠃$Yk2Ov��T3�jYZ^�c�Ī$�H�V}��n+N�]��UC.l��	e�ŁJd�M[t��CYO����E��0d���}�nA�7_�Bء�xm����Q$X>�V��������Q��r�a{yba���[F���ۂF�i$�٢�D4|�8 W�p}v�S�(���=J�4�k}R��xՋӔ˚8������2���>��g7@ꬡS�X�O��;���'t�Z���	lu�@函��aEn3�g�X�-���Vu<��YT����~	2
����l\Bh�|ۛ�J�o8TQ�s^=JA�<g�]�[Z���S�N2��:+z
7�9�9�G �1��Cv�۫�H�j��u�$Q�Y��Q���Q�H��9����y��1���a���l�O�,��k�l/Z\��(=�-���=�!���Z�-���H�ԸG�s��>iL9�L��ǋ��\��0#A�n��1�\:�)�����I{��s�Pd{[���(�榞��o���ô����H�x���"*v!j�8@,$�԰i_����!��q5��5�Z#<��Vc�����%P�hՖ�l�N�t��-���~h�ܪ�k��1<��!,M</YU93��z�I��R<,�'�dx�"�<���.���U��n�q�MI�Z�~�L��η��緶��yK]�����q7�`�H�&e��<A�W��_~� yr4ڲ=���?�>l�7�ٸ��i��eؗO��ڎ����dj�! R��j�3�x֠�8�7Db��-([2�����j��`�Ϻ��e=�A���U$�9��Q��k]Lg��9�L 0"�����U�j��6�iq�ƈB��qN�e���5#e4 �m�%`C��%��پQ�F��ߥY�I:X��B�S9�	��V�kj���5OM<H!v>y�xB�m�!�ԫ�[Ǝ?��p�X��~o?6��R�DlOlT6n��U���
v���J��
}-��eë����'o�R��<I�u���Z���v�r]�H��߸��ƽr��g8�\�
d�L�󨴄�,u5j�A��	_�*!��y���Z���l���.z$�Ԣ�^�y�'3?%B�p!OJqDC�����n��Ț���"�*�2��'+�,;�Y�.�ի��u@q/��,��,�����Zݴ���_���;��+tI���{ۓ~Ҷ��jtq-�{6����T���=h9��6�:Aҭc��0���<��D�ȌbEi��4tQ~��%�`�	.�`Y6߀~0l�]��~�����ZkX9tߔ!!˰��1��Q:u�T��ӹ�ڼUJ��9�'�dr��N��X҃q��"����{�H9��w��ɻ~H�5{.�+��v�����m-�C-sE?��]���*\�3�9
Aaa�' '�_Lr]���[ـDA���iK}�:���2|\9�ڕ����ڄU��� ��f����t��.��Ғ���Z1<��GG��w�2��gp�~�Z�.cH~�����}�U�����lm�,�WX�g����_��Xk�g9rd�u0�ۿW�>/WE[�˱t�N_ݱX�B\����rݜ�d�؅x2�a�� �&G�1��t���BX�Ϙ�l�1��������I���\��Pw���MNbD"����n;qp��~<�Zo�`.�j�V�|��U0�?>7E�`(�'.���8"b�Oo�?*H	��6�.N!M��\^嗕� ,��{� ��NG�i:�ϩ=�p�q���d��r�kG9�_[��X*:ǀ뜊~@�#D'�Maqo`d��<z��x?¦�iȝ�r�n!匡}���.?��%��O�դ�a7}Jp���*��UN(���u��/�E�:Q�=\��r�0���@q۬�y1)"pZT��"���x2�0y��d���&�!1��{�����L	�R�X�Ȉ�0yd�t|~S7o��δ;�L�0�c#x
cpÌ[�LZ��k�P���	��"LfEK�^�1.�����5��ϙ%o-�iSoI��y�#1y��	q�x��+b'�����02&��;U��<�Ttgy����?^�;�a�y��;��~��$���Oo�/R/?�v�K�UDd�㋫}�H�KA[�˼/��1L�!4x��$��S��2XI۸�fA�F�I2�W��P@�b��o2����_��ih�tQ����TF�w��n���1T�B\���n��z�s������摦Ws)��	�Ҟb��:Hw�h���#ؖe�Pm���>��V3?L��������hLl�k�S��^k����'~��S���L'��W�=��~`3�
>q�mQ���@�b<�Jj@ϐj���6��/��dc/�<�r&�����ضK&��yh݌��"\��q��'* ����0M��f�"M}�z�k:�������`W÷�O��{��^~�ˌ�L�;+�6D��=~����ݓ�������M���!�����7��ɫ���~�t�L;��
�:�<���"��o�݌�!
�����H�l�nÃ[�\�ȹbh/}��J�U8����h�7���T
��3���'�ODf����k:��ʵK� ���Q� �]��Ǯ��_�R���	"���2�o��_-�6A�����>�&K˰p�x�k��NЛ�jw�J���$�S%~p�5�����b��vb�ctN�/+��c�>)x��u�z�(`x?o�49���{��Xꮣ��Y-���t��B1��w(��Y�8�q��Q�5:cY���'*��u�_��f�*Omo��������]'�4N�r��]G��@{�ڣD5�Wƹ2E��}Ls��v��V����d��6���6�E5@���T��9�\�I+RK���e�i���V�i���g�(Z8Y�1Jh��.[�<X�;�rn�I�Z��J��1rȝi4��z�=n�+cb�L	�����.�J��zϰ͓<,���:x������ĳ�ñ��,�:>�]� ����g��A�"�N!�S�j����u��;�	}eI�R��4�/���Қ�U�����1m;.�F\��L%�ɳ�uΎ��_Is\B�<H�&���8U�9�4����Q�P��Z�/P�$J�w�Ü�EmH��?�!V�Z���~z���R���E����9+�wt�vM�0���(!�³/���d�`B| x#vS��2���b
�<|�d������)a%�X��w ;ّ|���DmO�<{g;���?�>��Lx_�>��$<�с�ðtF�s�3��>��5x���0PȂ�h��S�Cα�o:jA�dJRu��粢T�c=�|�t��\�/�m92X}� �S8�n��Y�B\�N�Yo!I$̈����gc��1�R>���������H-UH��bѐ/�ꊆ��-(��c�+�u�����h��5HK����cڵ
���9�]���4�%	�Q��c_�v�_�ǩ��n�^(��� q±k��砨���<�����U1b�"D66s�� }ũ���n���\y��x��jW�eIǩD,�aXk�&�p�|<��T��t.��_�\�� P]o��x���n��j��g�����^{����)�h�V��} l�E�k�t[a� �#B��n�tOA��&bMr������`yW"������q�N��̫�>B�N�l��{�co�|s!GY"\8mu��ya�T#��*�ZMJ��
�
^�a<}2tZ�w;��˺o�[c0ز��9��R��/�����9a���y��)�>���Ŀ��nҫ���C	��~�aP�ש�]���,��H,�x�r�g�6'�G�f�T�r���Yz�zRj�G���5HW8/2�!3�	�vX��t����V.��qC~U1�Nrx���Z��� ���	~�Q���0�Lx��H�BTƾ��;:�?��%#��5����%�B�L��0�F��zp��-ط�R�6uXc���if���cܝ5���]S\5.༶&gr[���7�%��z�Aֈ&`����0�Jv��k\.����D��kp��!�G��5p=��>�`��0��t�"��ѓ��g9�㦻�Uɦb1��� Ep�f����8�i�V�����Β2p����x���q�C���'a7���<�9�Ǉ#�B�)j�2\�J�Ƥ,�E����ãS�I�jx���]�0P�U�x�<4�>'<zˎ��QY�}�1g�z[�S��r�#�����O+�pu���Z0��ɑ��q/��<����uN���۽�96���1,��M%�D3���j�$]��+���(a�a�p���@�ϱ�%���U�21��w��)�[��~�m(\A*��F�~���]jXk���兘�]�f�A>s<�J�)I4z��k���і�`�Pi�̗~.���>cy!�����\Ȣ��*������pvm��0���<� ٢%=���tFЮ�އ)Iz���K�S
t�����{{�C��~	�<�}B>�'(f�ft�s	�e�A/���3�	�{�̖�i�BX�>����'el��p�јLOa��a~�b���&=Xh� ,/\��o`xHaf����'V(a�e#u��	sw�F�V7�����E�4;h�~t�f�b~�/r�}�Pk���Vڊ�s�C"\4d;�W)�oZ��|8��=�Q�MEq��%S(���#�\l�1\�l@��"pJ]�\oPz(��OqYj�7���wm	}�nNW�Pp��{|(�C����.�iC��!j�c�	c�aAZ�Hq�Lc��z���\�k5�]��5.�.�h?�TGt��)=���y�ң���S`-�V�����"��{���I4� Է�SSIm�7��uа�-ҋz�?�։���K3l�fa.K�nEo�.$3�PvE1c2���ɏ�]n�����{� ���
}�o욥m��V*JQ+���Cf37�o��d!61D^Cdj+]>+�#d5���&S�ulI����Ɵr���##��x�O3�u�HP�OSo7hz������ �R�1�n&��1��/�X}�	4��hg8���Ȕd�����@q�*��:�)���rɸF� ҷ:��q�2=�7�X���>l����:��G�%w�߭~i��c1AeS#N��u��#�s�Ѝ��>���ˏ4G�qc������V�qlxl��\Mԑ�x�.����j*��iõ8�j���!xE��k\4kݜ��~������㪯�V��nw�{���C�Tvw�
��{U���z� ��&�يTqq���5�W�h�Pc ��zV�q���y�!2��� =d]�Dޔ�{��_��hi��\Y����κ]�tX����`��#�0���N�a���?0�Kw��W��369�'/�lF��Ӣ��
���m߽����]�����:�|P%�o�>bx��I 1b: �sΆ�+^G���c����" �L>oj����6 ݺ�"�r�~A�=>d��s �֘����N�0��䇋?UЍ�V�&���=�Ji��}Z��	Cv�F"����>e�[�:28�&��Z�c��կ�,�y��|��ÌK��w<~���7	GJ��֏�.ݥk�LPhm-z)6�~�T�I�
��N��~*x����ӥ�wܵ��l�\m��\�a(j��Q��lP�;#-��vv��}Ԅ�[��!K_���`��v�A���Hg�H4��gG"���'��1]ֿm��"���T��M��5Q��k�ɩ��Gl_���k������2~Ԟ�MM��)-��M7�����S"�%�i[������d��u�Pl8$_��盄-DX�:�3��}9����]�˝���X�ۡ�W�<�}�63V�?���+�I��U�񲱪�䅿4��u��" ����v���+&[�~��
d*_���L4!�`z�er{NKb�롡�{�!�Y����j??$	$���Ԟ��6N�[�$P��4I8ˎ���.��(�7wG��B�����Il�8�{;��N��P/GÍcg�Nإ,�Pק�\͜n��jĜ�@s��� ���J|:��EN��xAC�ᔝ_Z�8+��G�Ɣ���}�J7��;��o�h��&e��7X��Yufxjx
W��Cˏ��>>锋�¨�qH�E�
F��-�w�N]c������I����+�#+�_�yh�Xo`�u�u��"����Q�ۥ��?�I��0+:���=���}���X����Աm�Y�>n��'�����ΞJ���e�ץ�Q/��� ����:k�"۠-�"F�s*�=,�qS�x»b��T
��������.-��)}�4��Lq��6�5����heo��@��\S�e�����d��^�,:� l#nk����kS��}�WД��{T%�Ԯ�Y05s��y�^&!��Dh�t���9߄���۽�Z%�{�s�/)0�2'i��݇f���U�tB`���|�fڌ�-k�[ˡ��U[=���M��g&�J0é}�����sl�?&�4I�PFM�z/�P��]�5Ҧaf7(�4�_��J��f�� �`��s��J<�BsY�$v��鉷U�ƩC�P0N3`fJ�N��[�bŭW�݆L��*����ی�#�u�lcN ��K|���03�1 ڲrk�[�N�����Pz���[#θ�O��Y-h���=����'ͬ6U�v�р��7y{������(��M-_�6tA_����)�GR'�0�땠or�֠�dFtf���#������c�ak�!���m��ڃ�d�����1��J�ھd�\��[.��@�{��������u]�q����Q��t�`���pw4#M��0��L]�zdw!%)O���%7�Ӻ&����RW��Ŝ�aj��SѮ:惥�A\Q�S��ǂ�G:����,�����Fl�-���p'�'�fX���D�}��(Lo�WK�U/�J9�S�C�}d�]|
|5���a��;���&��C����M�N�IT>�9,�P����g�r]�b�js�����½L��Dh,h�]���2�U"��W{"�����'���?vguH��[���p��&s����U��Y��ɷ�,��B��	f0q�4|������ζDڤ����#�'!�	��TV��=
U�߆�N�ٵ�!�������i�<+Z{���h��T�z����E<y��X!]�^���/<\�d\�K\��}�C�=_G��a������c��ʌe��z����r�2y
	��,c�U*�.�8������Ǎa�QI����U`����xܛg� f\���׳&�{4i�oSZ�[T�v���2R���?/���R�m_�׊H�G��b8s����,�p�D�cpT��\�r�����)G�n������s�i󿮡�Q�	���+z�fO`ID�|��n�@�����.1Z2��r+�^=vXAj�V@e#u�_� +���E�+�S���$DB�ʩ>��>����i�w-'�dwBz��-BP��gaA|�0ʢe��"��:�?�@�"o����z���c~��+���]ݼ���9v���+k�[��y;���P��|9�f��C�B� =���T<&{mv�eL,CX��3@��c;��/gΨ8ym�hGr�Ն��+V=�浀�,��B�+��_J�����?վ���B�(�B�Z�d�&����o;Q���*��e���9����z�+�j�D�%��V,���W�؟j˫l���ZfJ���5h������ıi54�'H.8��%X��b���&����ekE��U:�G�&8�[������L~l��c#x�O����`j�DyB�w1%��_G�j�X��9�>Qx)XJ'�3�[| ��
�h�m����76�U �˪�,��Q����a=}�\�t�&�7�Z����k�Oǌ��69z��������A���x^�d1��R�G p9y9��< �t���.��|����=�K�Kq���!�^k����i���R80�;`��%`�{
_�S��Xo|�����	���=���]/NTE��!]�cK#d��l��T��5�\/<���q��'?W,h$��O�J��p���O+(�8� |�/K�d9�E=0��-R����0n�(1n? �j�ه�e.�T�׍�u|�4�-F^Me�P�����jUI$i/Յ��qx���7�lHҋn+��!s���������T�>@`��5A�h=wS��a��&��w�I_ì7��yk�fav��gZ@���F�Ӝ���Y �]=l���8��_�vӊ ���ED�Bg-�8�y�:�?�6���ͱ�ܨ�>n�����q�ݢ�5��R�5��?�X��p|�R�
�RK�ǀ����fV�7���.�<ή=�����a��R�5�Q����%p~:u��ߋ��]R�u�8�r��YA����r$1�f��D^i��Gzk��)����ސ��^��J��ZI��0��� 'q����H뺼d;�6��\�	�QWL�RQ*�Hle�Β5[N�qqr�ܨ�#�"�[�ղ�[C�&�[��t��F�P����@�h�g��z�%'1�ΒmJi�q��t�$��Ӡ��r���P2��b��R�"J�p������:�>
��E���)����~�N���oN�x��R�7v�94&��Y�����K�	�E�S�.(����2�t9�6󕷚$� :��Iڮ��w�)ض7��^�'�G�l�#5�SQ�*6�r2�R^H��z�`���$*`M7�u�A���M�@_�☚c�^R̈́��6-fnL�$�u�6ޞ�_6؜����Fq��9xv�௣f�nc�x�OsP.*A�=�D��ί+���3�ʋoOV����+��h�"�8��R�r6X�I�\$'�i�q�Tz�6�������fQ��yą��o������~�s��ǎ��D��E�c|9۰e\���KBl\�i�W\�g�@>���5��t�����4m (���@���ҬO�Y�����#?Nu����� [y(n�b��4�������6���)�h�tz�
��U�խ�2�z��Ԗ��"�m��'�׮X���I��A���c���&��L����|��Z�^��K}M�(��R�%'��H*��H|Z	��cV��Ё�&��!�G��t�[�3��d3��ո]Ě����������i���QKu�Y��j4��캢��ICǿp���\�\��Iw�9��D]Z䭫��om5$�LAa6���z�&�ީ�ׁPc[%�ɖQ`��uϴ�a����Ek����Q�9��FY$���R~��e�
�Q�9�4���T'ǬXǹ+䣠H7��r�I���aJ�#�D�G҆���(���@��e��R_��'NY��;�����>��`��S��N�Ąhk�4 q�룿VI�_\Ǎ�bAnoa������4�#M�)�Op�8�0uF��7`Gb{l�$���E�ܖ��B⭙!�X];�<�DFLz��Y۔�ߎ���ل/f�ƹf����������N}�ls��KrT����GRS*b�rYk)"�CNf� Q�
�PyyӴ�����������uԭk�j���;�&�Z��̢�>kK��EU������򗊩�R�Lʋ�8,i2WNx���������C?�Mh���۪MÜ�lKZ��L�قĆw1����a���5�Q�o!{���wlk��;#O3�5�l��T�Xв�Yg��,f9�9�J��s��فU!�?Bq��u��d@-���&�Q!1l���t�	�c4W��9��T���s׺������U]:��G��̿��c�1 &q��E>Z��Np�qFL���-������E��t�'��Z�}�+�����Z�-��Ip8���� =���n&��ћ�c|�֞�O�1狿b�M,��\I����7��.@"nir����&�s�`���C���Ƴ$1�DPqr��}�%^�UWߎ[���k8��4$xaT����nz+Un����y���g
 ��K�ˊ�Ο����!:)�܎n��h13��r�[��4��ܐ	�eO��i�L�T�PY�`4����~_O��,W�}�����Ъ7�Etܝ���T�5~gB�d
��*B��̽�0�6	|U�k�[mg�8a��u�N��_�]�7=�>�5��)���3{b����C�~H)1�u����Q�1�{�e4i0�rp���f�4Ԉ*�����g��
GW��+9S��PaH�Cn�����{D3L!�A2�O\悄.2��2�c��N3�}�u૑�|3L� U�KB.,Uc�r1v��}�����{��w*O�����z����J�Og6;+�]j	.����^sA���&�9}=P3�x�3,��� 9��Աs�ʸ䈯{�.�Id�2�F���8;�� ֕�i���$J�3�L�H�5�Ga��~F(�c�ʩ�zZ�����?����;��ۼk(*cKO����9�����)e�P_�+��^)fD�{��T9����p��O�G�"��P[�+�v��UCy��X�%܋�J%��f ��Bq��V���eN'z.{_��ǇC;o�?E ��<I~��wWc�Z��dN��;%�V>{v���E\����$\��|qi��p��u���|ǹ�CLh�����5����Q,T��`�x���RI���|��������A��|=e���Ą~�G�i�m����T��X��;t�V��	�B�x#�'��~�&t�#b^��D�������P�M���#	O]*0�0�%�H�B�V���tqAA�SX�9#@��$\�6���ӄ=��b�':ח�#�Q�w��rF;�r#�?��ެ!���R��B ��K�K�	n��A�իzC{��@�8*F��7F��b����p��\� �-|�צ�<�)������렳�B�қ0�9���hz�3�e��nA������l�M�,/q�0�"����z���~������6�����?1Ufa~ o�I�J-Auj��4�/ß��̼5�����,��������	�S���X�73���l#��a;x�:���A�����e�:����[XfMޢ�H�������.��;�aB�~8[K}�����I�{ �ДMy��U���%|���MFn]�,�#��c�תI�X��\�6}�������y�N �"?#C��'�a���e�kne^ݿ�׉�cP�Dē39� P��ܡ?�4i乪������g�#��^9���lH�e��v�rx/��߉q�~�%+L	n�:U�q� :62�Gy��@��^fKR-��(���( @�Д���8�&��.��F�־Cx	5!�����?ξF��L��{s|=m���}K�4vL�yP�^��~ң��-�/#v����:o �ؼ��xO�.k�u�x�'�XWRB��b��!��G�xi|�3ַ��*���p`��C�	T�Hp�bM,*bB�P����W 7(�X�ѵ�&86�R�C�j_�Y.�[���W�T)t�ƫ`��4[��{؍Q�G���ǘ`�	�S �i�-��m����]�f���c�f�z��P���ҍ�J\, ����ȑ�!ț	�{_��]";� h�(����@��{�s@:@�H7��w�dLu�g�hY�!�5I�k�#�1��5&W��+�ˠ��	ܭ �����!��Yu�O���>�vt�d_�b��~2hN���Ҫ%i�~Ƞ�u��o$�+�ұl
�H-˥#K�r�h������t�Y}�O|m��vW�,��_�U�ۥ��O�姐�܏�Y��Q%���h�zQz����R��_�����]������#�|��OFQ�#� gJ�u�~��<o�[�?>�x�A|u��|*����
)�c��B+� F���#��{����Z�ͥ?�F�Jx3;�$��!���Χ�}^%�%P �����tm�(�#�h¨$l�0��KjF�y�<Cޘ�E�	�G̵~���r��RBz�ݶ���B��Q3��SNO�4?��UP�s����"��q�P.�쳕.����?�x�@��P�ɏ�&�D�|��ذB����szO�!��Ho}`{Z�ϫ��b@����_Y+���\f��`�!1�u���*$O����8аh���O��)3�H��X3%��R$�Z�!���wb����/t�����i}��Q�Ź7�xI��9��)�����s�D���1Z�1,���-<?q���A:m�^��T=b�"&�y3�|xTtÇ�z�y����mO��jOġ�����L�@�����)
�}_�a�X2*��
�ށ�� ��2�� ����8���P��ޟp���W�Y6�l��5Mw��q0,������t�b����&~k�;]0F�Vzz�Z�@Jbf��t�i����؜*�.�o�(�gv1�'��HF|]MQ�Yj}�T����bwj=�S�-ܑ�-5D)k��#RB	�Ԉ���R(�ϼ�᫈��ΚOX�M�=��5|�Uz�Ԇ̼`�r,k�(�U�U����St]��0PNU�i'���Y=m�jY��+Q�_����������"�*;��
\��^M����5��%?��JN�������O�\�~^�ta�����1��[�X�.x1���/*����x
�y3�8s�P��jݾo��
]��Z���l�Z��Vk����R�f�����']}J�͏��'6˝�'��{mH�@�}M@P�b�$�l�~�����A�L��2��3߇3;�96�x�&;�k�a��mH2�S�Zb�Jf6��jm�w�G��Y!?k�e<��;�A���;�CR�b��SP�V<��2��ݝ�
�=��Z�~��Z�G 8��zef�힅�X�q�g�2����`�՜�H���g�hH� ����p�������G����ФN�%G~j����<�d"PS�2��<��^�β��]��>V�<	t^�%TR�CX�����(�Ѝ�P��:��Bj2��&qq��ӞpUWOY������$�{�o�U1T��9����2j������;G��/.Fs�~C	��A�/�ᦷ����R}�P1k:5�+)VnB��$�=�g�����b7ϵ�p�(z�
�������]��ͤf���K�Le�4�?(�A���Q [c�[x�q�u^T�Rqc��|�2'_��g�T���ʩ(�!��Wڼ�l%#�*����ϒ��j�G���vp0ԃx-lB���I�O���m���P_�&����c��e�衸�Q�7 ��}M�B��-� ���#?o��T<��dP��3J㞕ކC��W�-�Q!�l�f4�)�;����PZ�6��U5`\��M�K0/�;���K%k--���F-�|G4<�� ��ء��^*������,�[�#I�����i�J,�V֋�C9��J]�a��I8������EH��T�WƄ��+���&��ͯ���F�%���L3�U.�1���g(�{�ø�e 9Y��xp�����á�ɂ9`)�A9x�-�>�:�_��" �Q��4���qIw�nA����Ohɟ�����PN���?�]�1CĢ��uctO����ы'F�����4��07�t{>��~�{|17}Ǣ���]�*&$*�OSz�1����E��v� 3��>�E�坧MA�CZ�6�~qg;H�Z���,
��~�b3X)��Stwy��Lj(w{��w��u9�>�TNK�Ph��Xhw�eX¯Q��Уoʑ�䵗��kH�����r:g!�$(��8����7D.�M}�\��@S����9/Gl݇H����K�|�-r����Fʸ�łB?C�u9�>3>�,�����v��n$��N!�1p>%���b�arE��y�� 3
?&ĳ����PZ���Bh�Ni�Ў�oUDhT�D�B쟱
5f��H�=b2/���ᗹ�t��
��B&�h�-�@�;,k����uq%p�ԋ=(od�g0tŠ��jb�>[i~�s�kben��(9�Q��<��aXYm�H��Mz�tK�t�$�
3��Ls������\�B\�9%8��G���`\��<�e���k� 3_����TGZ5��.���;����zjk������[�ˠrM����]B���=T=O/�#��3"
c�{���-�؀��4f뵝$K�~������Z�%4g�女n=J� �=��f4�{�_X��HxCwe�O�I���DNg�3��ѽ)�5	T}��h�#?/�-�t�֔j����ԎY�Mlsd�?.��$n��������7�"�G0܋�=�o��_ �����e�ܶ�nLe����\�u�b|��	�MH�Aj�٠��Ox�����#����f�H�H���yzV�,3�Ll�k}���ڼA�D�T7�*Q����#f���� @$�sq���m�pAN������5<�q�}��F�楑��x�P�?��_�8�|Nm�Ze��<ѷ,�k��F@�Ay�V�3��)���u^�w�m�&L�K�­v�r�w
�ȹ�P�\"������/V	޺q�)�r,�kBK[�J����g{�Y�$�=��4;�=Lh�ƈcЅ@�x�^�I�y��������"ED�]+��.���&��m��r!�
�X�s�V��<n�N���;cp���냨���G�k�Է�t7�8!u�8���P�f�x�ٻw֑�*�?K�@�-}�|�_c��f����vv����h��xX�{��:�����beFN_w@��Px��Dfi��� ATOÞ��k��e�����<��HQ�+�9�u"W���(�@A|�i���ma���	X���˷�L�wiw��iE]�����0ECW7���l]%����~�#߽�����t��n(�f/N
>KA�B2#��6��$Y��0��1�'1�z�߻�t蠷3�e�	��Hz���y������LB�r}�@�n�'��S {�����X-1eέ�a3�V,m�4~�����#f��C7;6}#�'_"�D�;4�f��)3�t����G�Y$�!�Up�z���^���߰�/~�������t)Y����M	O8&X1���-��axAE��bb$B�<V��{&z�9��9���3�c���X�����ۿ0����o��|�r$[�i<L>��4w�V�j۹/U�/�=Hՠb����m8������W�>�V(�vQ�#�9؄H��8黛8|u���8�)�,��9{+���q���\><��a����%E"�GUA\3� �~���0p�<�������/�a�3���$������WPO�ޖظ���I5�·�N�Zo<Ơ��)�3�j��$L_��Y�أʶb�Ob�`j��c������t�%��o�����a��va��0֧���I�]�h��:�}$�u���-��Oz$�ڪD��6 m�}�,�/�V݈ʩ���	��a,I���,���X�_�D^C��y�V+����ñ�:���TS#�s��F9E�2������ٽ�� f����́�;1pG��"��&Y��+bK��ZJ�|�\�lQt/"�����5��.��0z��� cE�N�A��g�B�ћB��'}����"0MQ�8i�D�Lg�@^ϼ����p[����=S����̼t6�
t��Q�T�������G�N]ZaG�\.�yu����si�H�%�)��h�m(�\֯��9��I�_ s(��'�:�5X�X��kfhѥ�r�6�b����ob��¢�O�pP
��% ������ռ�t��̊Qޮ�'��w�K��C<Eφ�O>A&<���[�>m)�]�=0{����� �wV�ѐ@%N+KP"�����]@>=��jN��K�MxbҊ%D\?S�t�q�d�hq���,��і0����o���%�6�t�O��e`'Es��&�5m|D �P7�f|�aP	�v��(�.3T�w�S�"�b���B��(o&=+�f���c�Ɵ�r��_������~돇��A9��䶰�p�ޮ��Q����1(���;��w��H�9�&JF�Z����6�Od�UY��'[O!70�f_y��
��Ve�j�B��� �~>;=.���f��*d%�4p��!��w涱>N�&?���۝}�a��񙖄6��Y'�� G��I�G��ѵ��eP�T�i��_[�S��:�%�t�6�ˍQ��tA E�3��r������^0�(Wu�C��V�/F6��%d�J?'5��؆8l>�ף���U����y"c-CU�{��7'�I����(p��� Oq��aI�}�+��il�3_�
n����^-|p|o��P�J�n.j,\��bۛ�ls��E�}<�SKB�o�E$8ܓ��QCBE�9)A#��+8f����9Ͽa�4ݼs��F����ͤ�g�*3�J�� v�2z�%~�shMdj� �[�J��������.�a��r9x��X��NO*��w�W��b���g'Mҍ!��5ȥFL��z2�/����0�a��T��/$U���F��n�GL�-�Prq-dbT���,P�1����T�⬹��4 b�3���䐠��[S�	��%|y��4F����Z�12`L�ݍ���E=
���K�i;���
���JL!l�F���E6e�����
k??�AL�UN7��'���ˏ
Z��f��q����\�_�0bĕ��Gh�@�_����t#�{��	Oag�2Ȇ��A�P��Y��1:�	H<o]a&��e���Ej�:Tt���'��"��cQ�A�������ۺ\:�m�CPd45Ե�]��#K0P�`�������9�DӁ��хf� _JBtj�Y&�-�uo�M�qLY���B{a���V�O1FU���.;�;�e�޿��l�%��4�zϼzE��� ���p>��a]Pqb�.�|�UR����Z,2��H��0f��F'�w��0��6t�:XG�
��hz��@@�)Npa������o��ˁD��Ԣi��E��[ހ� 3Z�����=7��"�)vC��,����xh���PDQ�cY)�E��V�(Z�D>�F���~4����ث�ӭ�<�M�X��C��uO,	�ݚH�U�`�J�0/F�Z$��Dx��t�du�d�2�V��HD��z�t[�=�"()���`�[3NӾ�)��?S���z��=�v�r�(�丣K'�vS���
�Ƞ��okd���	4��Mƴ�|_j��몛ڢ��.���������Gkm<	jo����k/�.�kR�еF5���f�Ba�ۅ��d��~��y�����%��z���w������)ܢ��=����g�Y1��ˑ'.L|��V�EG�/V�Pe Z���4�����MM>�|E�rL+���;��?����q��~+vR����5rQ�r��s���"(�ҹ�y�z(2��C��H]KVA2��S�|�H#v����b�0F��L7����C��2g�D����x(��g_��PxZE�H<ɖ|w�a��W@zۀ��ba�$s{l�Se����<�Ը-��κ����w6��~Zߡ �
���Q<X��@���XO��`�irp����<$��dFY-f��Gm&��f�#2��`
&_��2!�
jx팿�sa��o��@���0�7��i)T�H�W^�Pd�Y���4�
<ET�����M���x�@�d����/�{"1
U��B"��J��H@8��⹔2:�S���l';�C�I��f��e*bx��Y�	�L��yO���c=6��x�َV�4L:�.8O��]Du����R���"k�1y�z���NEa+҇�G��^�Dw�Xq;�e�Q"��R.�������>�w���w�[��AoQR ?�"����ȓ����	�w=Q�@?�|��+�Ḁ����RV���kl����zk��%�V�QX�Kp��J;a�(jX�&:��ʾo���������T�z��}k��~1���b�I�1���pן]�&4�Zn/p����fb$�&&�?�O�x^���=���}Y	9߸[��C�g�*��'Ǻ�r0Pu��arn��?oV�{
�7b��n�]�IG��%�[�qؙq�u(("T���o-�`+�,8������$��LS�?N��x�$;���D�e*�Y���C��X!6�w�`�	*�Pܟw��:V�Ү²ϡ�	bb�}�}����!�٘��&���!����5I�ԉ�(��|�/k��5���l��� �=>H���ܕoG���RpB5�wMZ�[ۡ���4���	�M� �nB0�}P���4��M�_O�j#0�uH���	�1� �Ka�a�V�\�P1��"W�0�su�/}-9�\a�;f�.���:<g �V�>���J�������R��_C�I.��̈�>�ա֘�m��^v�r�hB�R� ��
m����5��VP�Vԅ������RW,ہ�}�2z����.&^"�] �ͽ�@ �3���;�N���D�c���Flp��Em0G]-"� }����K�֬^j�t��e��"�S�b	m݊�f5"�	`�fQX,�\s����O����u�B���Lc���X_��\���̬�^ɾ$�}����][�(Q�ml�F��1@n�4�^6aԝ��O܆.���@c�W�\�U]�9�Q{����/5_�3c�=�OԩG�d2�!����ԑ-�D�p��P��NO􊨟��`R���ȓ7�"W�|�"4ϖ�]���hp�f��Vi5<��9�|���j�va�R�����%���ÝN �O��W<<;�N��U�C"�E��p�?X<��g�ԭ��Yj�;��H�b��=���Hdfo`9ܸ��$9�U�PÏ��I�c��;�����ru/75%��v�FU���R�5W�K ��roFs�Tб4?�U�|Ӷ~3�����8�J�jG[e�Ryܸ���3�fà�}ay*4�ّ�����/�g�fy ���T�W1}~Wʚ�v�  D�: G�{�&Yxp<wm9�AHh�o��@�P��r�+�v��a�:�Z�@�s�n�tnٗ�4��崜7c"�u�WB)��M��:�m�\�R�6�=�/��"W<�9�ΏAE*C�|L�>�n05`�}�D��D��R%��.Ƭ�s�Md�s��^�)���8"�T�<��ᤲUmw0��v�g��f������s*�N*mu?��u�r��@)��9\BL��q�s�2�F�8������0�U˔W1gu֪��T��Y3a7�uE���*��h��Mfy#}P�2��?��>"=�C��d�.��_��?���'*=c%9a)�9��,x�`����l��:��6q7��"���������� _�K.���Ux{x�zG�3�-�	��;|o�Q#��cKn&|A��x9�bS}���@;>%ʈy�,�
L��h�U����t '�Ds�@S�yN�@���B���[� Sn�g�$�b�yt�(^*(����ɽ� ξV_�p����Y$@����t�?�:_��sm]h4K��'�c��/��
f� ����a��H%�g��N�+�u{*�5��v���hJ��a�ϩ�<�r�J��f0Z�p'�+�p}� ���i�b����Den`|#'T�dюe�c��݊'5��&����#�Fr����=3��8�ńV�{����,ى�h|�K=�F�)S���9�k@t����)�	 lsy�GO�n\s�2�pҲTw�1nФF����35J�v:7(�'��N�a�۱�U�ط����N�cJ��M`-��DW]���M�@��y��dʬ2���/QV�|��ݻh%���$���^8��E'�(6�!������=�T���v��A��]z�s�K 1�]+��[�G͆���}U�Y�	�Tm-4��re�
�����9���s&s73J����
pP��(p�7�1��s��0�}�a�>� `��t�K�.[lR�#�W�z���:ր�̆��p��Q�����J�t�m'�O�� cefL�n��]O~�����L�&�Sc�U�I�R�O���2�Mj����l`�Sx3�
Y��T�j�Ko��/N�G>l{��p�m_�m7�1��
�{j��8v��o�݋���!�b�B�*�u�M[����)�-ț0��*�P��v� !Nb�~�����}+���w� BN����
���3<�W_�%d�~@f�	��]�CY��8��ϓX�ط���0$Gn���uO:7$,��М �w��էtL�Ne�K�z��>z�ewR��Q�)�b���?����gz>���؍��J[�3�krͤ�m"h��o�'���!9y��ܑ���������:��1m U�.z;K�k�������`�⥍nTrk�f�B��q���as,n�2&牑3ʀ-6��H3����sU�:Q�׀A̏��D�����:۫B����q+�ď�{�N�^����#X���Rm[Jn��^��B�{Q�.�ԥ,�� �o�s0��}�+b �:L�hVc��0%!�K�9��l��y'�yp<n��J�E{c�<�#��,��_�:�ޝb8�[����Wws��e9����-�Y����J�ʸ�y�Ym��@X�A�9K�����F%u
��o�C�Nz!�(�vGb�4B�ĖzX��&���?F���d�cH ��{0�m1�t4����!���#��f���+�v��
B�&ߗ:Ɋ��a���)��Ѣ>*�,cc>�L� ���-[��$���2�~�gb��x�6���f�/S�K����f,&��Y>A���g��B��yn�ǁU���_6if���#��H[��������7pU� .g�+�z���,k��]zδR��9�#͒vµ)��f��=NS���"�ZnI�Cݽ�ہ�s�?e��2�) �z���k+;E�jg�-����$a���W�@M��ɯӺb175��������7:x?����깶�L����a�Ԓ�%;�@ֈܩ�\h5�k���o���x�D	U2��y\7�~�� [qHu�dz2Za@�����y"����w�jhaǲ(&�Ġ��y<dw������u��v��D�)p�՛�2�-a��:�����������XE;�T��ov}ч�^�Y�}�nv?���77""����-�H[�)dx���0��Z�g�S��hy��Q�46�����x��/���0�-ٙ�+��"�J�d8�A���uG�Q�F`��X��|��*כb���|lY�$����jަۤ���/ ��x��0�6��A���s#���Xn���g=l�T�_
������ ��5��C�
O�8���K��C
�:S���m+	M�ۏS��B[ϜM�����ѫ7�@��l���xH1��zv��/�%{�������K���P���/��^���.6��N�X�����t�{ w�����ju���*��q}ql��.����JRk����8E�*5O���;{�/�Oq�����ieT7o\��_.S��=��rJ��De7&N���/�W9R)[����S�������3H y
�Z������ ~�݄ٚM��6kꊂN �0��t}U���+�~,'c/���OTX����Xw�{NZ���+&m��ltm�b�4b(2��nħ/�dd�W��<<Q,}�<�a.�3�����k(�]��ao�I��J�~�wfR6���Y"���s�D߶x�dQ[��Ce��<v7�m�3`�����)Ԋ�u��ĸ�g�.��}��o1u���t�F� �7�f��xxӉ�Ї��j�mx���'�����i�T�'��aJu��œ5�.��wV��I�,���O��5��-��8A�=���2WC�W03w���Ϙǲ+��,%H��A�G]9�?}8]B�}�ɯ������j���(Q�ʼ��=`�	��h*,�b�I{��ܣ�({�#5�13\����<�������"0sI; ��i�o8�TNX=[��?�����>ԁ�����Q�� UxnV��yq�����
v��]�7��蛰�����>��}���Eͮ��'�M��Y����;���l�o�Z�\�L
���P_�J�i����x�l���F�=���s�C@��.��^�0��X���pv�*�<5����p����K���ݑ�v(�PV?�6��rp
�`�-g�SS�*&o�Y��S������3�yf%u[���ҧ���W����fG�}��([fe���36��}�������R�%Կ�l!��{@�hN�1?��oϰt}zC7G�GtRuWo���g�E�b!�#;���uPDČ:^�+�N�@�����9w�=+;��g�A�g�r��Ǧbs����xl�w�o�w�O万�3�P9�;5z/6D��t��g֢���-��i�At��,�ǁKs�7��Q���7^1?���1~p��x�Mzt�}K���Arc�6�9U�2��{�ʛ��nK�a3�����|U�y{���/��l��CӴK3��(n�{��|E���P"1pZkB,J����z8p�%�������O�[.^�J�T\�zc�����Zs籴d�:�9�,�V[Up��}9����:�C����d�P���t�*vPP`ba�&R�&�*��)��}4~
�́�b�	���6sww�g]b�w��7�r:�ëJՈK�uJ���{QY<�Rf�J�I��c��6��>ω�:-��I!0��g��ӐS~��x"yP~��7F.ɉ���k�%;��v�MOn]��� uKŉ����]�͛��ndO���vM�M��@���ir��e���?����Հ�.�yqa��|ߚ� $��	T�TIC9<���G�uj��"KG��n7j��Rt5��m�#f![���Lʲ�JF�,QB� z��3G���ڱ����"�g[�o7���=����W�4��x��z�B�|~jLi�]�4Sq̃!��Iy�W=#���3|�c��R��V��{s�5c�H����� q"�&��A0���ϰ`��(��L7Ii�
��@�é:P���o�458 �
����J3�G�p�8IG�#�*�;�l}�ǀ�দ����i®�5��)�Km2�0�Ǒ�Gd���#���ñ��^���'���DGH�T3��Ly�͕� ��c�������3�]O���ى:����K��a}��Mpx�o
<�-�_�'��\9���lMW�_P ��o�9�r���4|?nq����3녂�28�� ���u��_a6A���Cm�b��R��:���hGm��8��,�.�#���Os���7O���R�$��I$]8YO�a�X���|��&�R_<�L���н�����]�v��V�����J���$�حS�)q�O_u�����&��:�r,8�V���7��,����d�G���5�gb��pQl����H&H����6�/,�1R��G�S~_� 8�[����E*�$m�J	��\1U�48�m���
�����X�ޫ��|Qv�sr.�#�L��P\u�r�/m��P<FxPE[��q��}{	�̴0���� ��ʓ	3����*�4�U�r��6I��F���Z��mdS��a��O���\*V���bK���>�#��u�[�Ü��7���N�UUu`�m�2���qf�f,�`K�A������<Zh�Z�ns|ǖ2��	�o������Xo�����؁�?[ne#QX#_�O��ܯn] �=�������n�ɛ渋p�Oba#$���,�}ޠ�����\�����}����m>�M:qZ#M��(j��?Hף��ϱn`��y�!E����W�B% ���*�_�$T~�<����`Z�|SKK��G,Ub�2�tj��7拁��D?�WUj<f��x��)�-��F���,���lOa<��ʖ��'ikk븷 P���X�0lU��~�E��ո{x�!�cc�JY�˄^òe��Fᴹgj��5���8�^�7�؈�o�R�j�(dd�d@�NE,�<��t��?�'�T�����	Q�7�Y�r����*>蟥ڮ�F2��Y<2J�jWB(�{�iW6��i
$��}��FWe� �씅����A�r~��}�RF��X��u�۴�F�4˙ĴB��򸂄��^PMu���A5UWD�꺸gd �Z�X�R0z�X��7j����ۗ_O����Ab���f�>O��J3�W�1Y2�����};�mCX��`N,3�n�DT�n���w��$����6�1C�Yrd<0yۢَ�@�����Vď��>�a�g��.�" �{'!�PF�#3��rF&*�5�`w�6���!�;��`0������ӈ��*L|eyg���6��7G�`�\��lВI~������2�y��ߡ3��oD���A�z�ԅǢ6�1��1�X;}�����h��i�}��?k �.��lw���h_�/ie}���$D��a�l����C�?>�|�uw��=��u9q�ŀM���{Bu���Y^}@E�Y6Xy}p�����n����^���	~^?%�����l�Y�e��:`����k��Agj�K�hZv���]�$1y.���Yqs�>/��t��xV����-�����Z�a�|a��6� �H�%J48U��.�ʮ��_��`x�μA����+Q�� B5��Y�Ҽz0V{P�z�����kŶ�ʇ��'����8�ǻ�O�
�u>����S���")mX$�0�t6he>�m�"p�[��
�*��1^ug��_�2��r��R31<�2����o~Q����_�4#�{P��Ԑ��Uyo�*-�@Lk�ɚ#q�8��� 臨h���7ߙ~�y�c\���6)��J���V�F��q.�)|����I��t,��uH��]6G��<�1�$iM��뚿��>��~X#������=�9�)���W��q��]z4EV@� �@{%\�`�g�KMb�x���	o_۲���;v�κ3_�<��}c��z��ڠ�$*�%~x�.L.^Ů17��|h��2��W��tĬ�����c�كBB�FlLy �!��o���щ��EK�X�P{{'�(�#��ў�����d�-(w�f-�zd��y�O!�?TM�O�+c��4�@N]����-$��h�iL�?��X�\COx�B�w�٫���������\	��z�尣�nbMEJ�?6C� 
,/�ݺ��Lo&<�yQ�ڽ�0@ƚ��:6sg)�r�f^!� �ڈh?���$:�C��EQ�⎦N���a���P6*6�j(`c���[5���"
�'Y��hd��Ê������	a��w�Ni�.�����2�̕�����v{(��A,Y�m�n6{Z}�y\1i����Qҳ�응/�<W����,j�\j'�qe���W�o��Z��g?�feVFu���"Bij-:J�ɋJp^_<��_T'���u�ɡ�Nڀ3Ńܨ{1�GH>v�w�'�IF��	��<���1RR�gf���J�GV��N�h.���
�2��0�Z���2~-�g8 ��Z�G��Wk�D]|��f���S�˸G�򫶾2�L:��BN�{mi��Cn�X�o�H}�E$��.;,.l��6ȳ-�W���L�64�ae3?�4�p�+4F�HγK%n���*78���I�8;�g�}5;�v��T��0�������:�c��b|�.��n� �2�"��|°j�h����5U�}�Z�tb�Zl�&�`��OZ A�8í����M|']�
��uQ������z���Y<]��Gq������9J����c�ruB�oD��]��R�ߚ�F��ໆl�<��V�9i[�����bʚ�0�A��.N�^����8Jb�4�<`�"�{��F���U��k���b�n-y3�Xv���j!p����Ƨ��y��-5Js��$��N���F��	��)�g00��م��uB����ޞ���7��RF|W�����<���,m����������U7�1�[�IvJ�mi�*o��`�p�&9��VX���u�IH5�#q����-2Z�$�a~`���}>W%�H��gN_Y�1�{m��qr��c�~U�x��l�r�[��g� n�`%(�S��e��@�|���¦>���П�@\�۸0κW	q�b;�	1�����1�lP�{��.���Z�r>,��ed:�_I��f�[-��*��ڃCmd��Y�C�F�Y�t|l��Œ�mAo�o����K$piű[���O�9c��pCJl�`(Z�nb_N���.�~�������E����;�Nl�լ��I���YA���L,�G��J�Z7'٧!X:)��G�kE�H�Z��SH딪�ȥ#*���.���i�/����;\3��鯖��稓k���I�p�sl?�1ϬXb.H��T�(�K��'}r�
#u�rK�0�,��^m�r\Fz��h0�?�v��t�=����f5���J`J�9"0���s}��+uIӝu�Q�F�T���nX(�B޼�� ���&�M���ƾ/Kc���P�'�K����\��f9mAX|��4c����~]<a�q��Y�j�%k/	 ��h�a˃.���R��"�-�V7���|��"�9Rёz�ۏ���itIۈ��;��ޘ#���I���[-Gf���<f?�'�1i�4�W\��ųR1`ѓc�6���go�Q�l�r�yE&$V�\Ĺ�û�h�&R�h%;a��M�54D�к��е�Ţ@�J���4�� 洮3�Z�~j~G�;���	9i�����`T�ed9$u�zҷ�Ki��hd$��7�S�(�ip�q}.'�Z���'f.�#�$�0v�.��k����߈] Ex��%�������;aA�4NH,ƚ\f(�嵐R{0}�I�7�����ަ\�n����Y����fP����c�=���һ��!�i�Q�xe��*9��֠�`{�S���u�0=�����d1���x��곸��9hzO�.M�o�a�q��V`t��Qp7-�d�%�{%�L�bF���=��P�({ـ��M�hT��-i� 'w��Y��L�xcb���4ن~�o0�#ǂǱ�9sd�Jі�ֺU6.vޔ��ܸ���#;�,������k"�M|�xk�/���8K��)Fq�;��I�wq�
�g��9�@��D��������Q�k�	�-�`�S�gs�Xm�H�{'DEE�߄�v�9�1+�Ũ��~�@�Y)��CO���c�D/�K\U��~�u�����l���"�Q(��/o�W�o�����Y�7��z"?�A*��]�@5�PJԙ"Q�#2Uox|3�<|SU�y�F��p����-&(p/Ξ�U�Rq�t+��ȪP]�I�G�O]N6�k[�x�y)�W�����M52��%T_|f�S��,ZԂ��L�jh��9z+�D�e�qY8�.ZGtB�ʉ�\�Iu������$����J[A�e�Kֵ�7���ܩ0؜�5L��ߗml�L�k
�ύ�
�h �|��Ž<�߷(4b a��E��6`�yn�	������n�Rn>���p�6����z7`�}JV�2W�V�!M����\[�<PK�V
��aD
��X�L��ee_ת�e���wkj>:��n0�䶋Ⓛ���E������XB�*U#a'�N��m��޲�8PA�ŷ"ϱ��覴}�2��e~F�tn�2�RQF�����3'��v��J�EwK�G�B�:�A��%j�^� �RgWFi���+٨d�d7�X�e�*�쫣0+���npB�&�yj���� M�0S��%f���=�'�K8�7|�QpJ���&>������Z�GfK�f�C/���ra>�4�L��r?�^a��Z!��(�W�	'�g�i��Ϧ/�m�lA���!��V�8����e�/d�ٵ#������إ�g���<����q�	�YSb��;�v�H����֤��P�~0��7ygo�+o�e�*��#�Z7���\��+o��g,��{�T+Z�0�S"&�mNjka%���/ݫ��Z��A�^������(W�A�r�
�����o~�?[���>J44>=�s_�Wre�]1|�jMgɟ�f���0���S	u�R|���(�N0޾y��>єy�1�ەɼ�fg�E>|���B�F���z�>?UI�%��+tl�>�v>��t���o��sY<�x< л�B�\�;��r�cn�]�X�oT��ȡ	[-���B���6���@����x9��
@��1��=��\���OX]�t�NV�	ix��lQZ���	�I������`����ۆ)@�F����NC~� O�Rb��,�M�AT��O#�qXR5�ܑ�f��ԗ�ң!�x�vE�8~s!�!��g��O��i�+�e"=FP��~(�.0�V;�RJH(��Y*Ǻ�U�z�0���AH�]�������Q��x��g+$)��U��Z��Bo>�GO��M�g{`�����Tz&}e�O��fxLU�����m����a��"u`�`_���`{$��X2+e��R���ַ�P+����+~��@�6�t[��,Yr�Uaw�'�KD �+�`�Qd�ab��Yv��o�s���~NE���Z0���/��JE'0����C�89JB^	]��d���i�Y "(�������aM|0t ����b^���~\���G�_�ހ���~�><K����ϥ��cc��������}Y�)�N`�&A�������+$hH�N��}�R��y|rT�x�5�j��;�e�}��������IΧ4uJ;�4��u�n��r)(E띣m ���b��Ul��JUm�����#���`���c(�ܺ�z�콄`S���{yq�:�����U���1���X"/�|l�v����g856{��vB��Z�^ٿ�z��i��τ�!�����^�oF��A�f3sc�]6'�����
v��[ps������ �Y�����Tڙ�j�^�/W�u(�	�������"* ����HWQI���bq�W{�����b���:�������'o�L�� e҇%7l8���{M_% %.��3��� ��O���r�L
Gh��Y$[��2F�|g� -���Z��r��w9{y��L��f�k�է9+R�.@B�,nW[�d؞+ k�aU����"�I�w�ߵU��>��~*� �E\�Đq}��Z��C��4Qo�}"��_}{W�Kܑe�M�/�%�O8�|:��
�l��޵'$_[�5,�7�S�� ���tp������P�Z��Pۮ9�-&,��f� �6��?�֍.朏�;���u(��W��w���ڰN:sϜ��}t��ۿ�,���nT�9�	�2��L�,#�[dP��X��iu,QoO�.k�}4���=�Z�ю��)m�N\.I���րY�	'�CL��찹�z�m����I+n�>S*�jC:��ᑊ	?@!�3��K���������?��hȩ|e��t&��_E���X�55eO��qWDv�&ݤd�r6'0Ƞ�����ze��FӖn�	���O,�J�c"��`HK�^��!���}��a���
-�������c�{�j"�Uf�d]%�Q���:5SX�C�������X%u�l]v���r��?�5~�ZFʲ@��v���M{V��"�Vÿ�m4l�����y�Oׅۓ�9�ܗs�Ռ��GF�y"B^����p{c�3x��~�D��P"��'���v�H���Kw��6��'�3_���<<KQ{�����bV8j�e�Q3簟2k��z�˂����Ym?՟hlT���~6���c=G�)�N>�Ɗ�R<a�QT�ވ���\z���]6p?�>��5�L�/!T�,�^H�l���D���Gl7�J��6��k𰚾Mnm����-��|�H�_5����-�:�.{̗p�$��{�P�&��j@�����Q�\8Q��AZ�Q�h�;�Nڬ���Nm��zEΗ����;�#�劒��p�zb�w���B,UlKkҤ�k��)��
�(�*�b��1o՝���J��Ј�6��܁;gg�>��n�_� ��f�m�/!�Z����������ˡl��Ng�_�_�33Y�-v:<�đX���b�fՔ��|ϱ#ҍ���]IRt�t,��5e�Im��V�=H�c�����V�mƈT���ڙ��ȴ���&�!%0�] D ��I
,���(���><Dm�q�q�5�ċH������SPn�R�-�,�TzqħY@�Iq�����^ �ƟIJ�>
��dY�i� �~���<)Ě�T�n���W�� p��:�aaZ�C���]: [� �	� u�� �iDm�I�5p�IeTr����ݒ����P��� ʉm鄭�'{_���� ė���X<�01�I��z��0B�wB�UG�-��s-E�n�P�J	��G�ڄ��I�� Ƞh?ewQ��֖�/�ᩢ]���"�^�kP�������P.ƶ��70� j�J����6I�!L�0��	2�v�I�a2�)�3����!��͹O3�>�ɹ�9�ܫ,�Uz�����3�c!X��F�h�����|�~=(A��H��j
�T��������ʋ;u�|�gU��y͒5ҀC/7-B_��o��C|��V�Ms���]K�B��A��Şk?�!����`}�u}������Y�4��bc�@c�ߐ��zRT�/�/T�(���I� �F!���z�X����w>���b1TIމ����1<���6H��jb���>=�"φ��gW�3m���w(�2�����1�Y˖T®$��!w�!�
�x����9H��謑��|�A��f����46��ޞ1��/�N�&���)�{XpS��8��,͸���	�@N�r��	�H��.Ř�P$�51����
:����{�Ů[`Gq��^����K�q�i�[{4 ���L ���B�ϩ�[�,ܺR!��
�H Y�x01Õ_/B�	2��!�J$Ж��˽�������I�ɮ$��ţ�I�;�F����<)��=��ӑ����H�3�\u�OĿ��!X�8	5�PW���I�$��9���?F;���]�eZ���-�Dw�hU��E �e�T)�$��3=�Q�x�{��vٮ�d�Pu�P�Uu.��p|v�sG��zuEY��$��M��Mu����&+~��
&�YY����������&����~p,�I�G�~`12�#m53��ޣ_����o��,(&.�+���x+��-��X���uH)?T����p-� �Gj��.���8��MSx�L�Q*K��k_*�z$f��cY�����k6��s���E�@��=X�
�J�����#��2��bMJR�k����R������N����D�dy��!^V���G,�;�I�mc��XP��5������㇧��<�,]��ə~���A�Hk*8?B�fo�[>��m;�j8�����܀5�����}D?�
5�"h������<^2;��=�1}�8��kU��9�D�Le��W�_�m����	��'G�g��������gF�8�����	�ڝ�"Ɏ݉����(�2���>&�X5��G�:�Z�O�AR�膖�iE�qKspI��k���ʉ��-w�R�#BqȲ.��^{����N��!�r���`�F#�h���6(�a�"��
 |*��-r��Ze&�R��/�����xH����a��5�n�,Db�'��gqeX=�|Kzu]$��֔�{-����@m���
t�r�>�sh3��٪�{h�g)�XZbS���p�����?SB���
_A3��t�y2��'dS��_�S�/��}��6&l4�����(J-�Pn�O1R�1�ٺ�F��{/ܥ�`�^s\15I����9]�)�Ë �}����������'yխ��%/�2����Ek�����hX5��I���Eb�� �+Ϧ��(m�U���*r��)�q�u���h�4�J�glTP�?�3�*&E���:����ZM4�lu�����z3��H��3"t��~�PLt>4唑~g="���P)��A�'ng3 >"��o����l�����u�Kޒ��^�<VF��W�o�%�S?쾇�U�(l�C��G��Ã\�=��i�D}�W�;T�8|t
��Q9̮k�)|�J�^*����7�v.X���CUl{TŁI^M�>����J�l�	%6U��[K��z`��	6�	TI$�ʎI��$��X^"q�6N�jKߠ�/�"EFv>%�8"���},��������Z��vq)�j���U�v,A��L�`�[O\�.R��.6���j�Q�W�Y1`YYs"�jS��Dƺ3�X���$��Aj�F�Lc�c"Q��6��i��A
oeFP7��O$��E,#���d"��M����Ӣ�Ʀ�# .����JJ%f�Q�3Z��µ�7���u�XZP���I�h?�14A�[�,p2�gE�{��ʢ�;���]T�յ��c��w��S�X������WY��el��$q~#�)!���"�/O"sð��1�͂��(�o��+�a?��i�h.L��"��5D9@�b��G�hF9:�{�1����of��i�}
 ;7B������ܝ�8�4�A3!{��.��|,�����_DG���0�>�r�z��@�l%8b�I/T���i���&b�5C�鈭��zǗ4E~z�h�i�y�nD�I�7b49��?�a��%ø���zco��!�y!d�KSbL���N5���\��H��(`!0y�l��_�V�8 ��W�x�n��mDksN�3#a��!�jK#ߩ���٭��m��޳�:��h	� },�t�P*,[������#��(�{%�CQ�v�O�ԛ��|6l;��(zf��#��Yja%ff���_已.up9�K�І�'{�R��k�o�ݹksp]�
�< �@�y��F'�X���>gud
67�a[���lP~A�&K��������>J[�*S���`~�9�qsj%���Q%�s!�>G-��ؖ�������#�E��2�n���d@?�o>FB�E�[D4֠L���-�?�V�3�s�@����S��q۔Vr;jx?�[R��ͮ�u�C�|�G�qm��+��ٞ�n�щ#a��d��?'r.:>s|��s@��zM�뫫� �S�E��.	����!��>H�:�B��J���]]Ó".���
a��vۃ}�gZs�''tq<��>0"�:^��w(~�b�!RC�t�@�3'���	�5���B��������^��NT8�(7=Ê8�p>C_L�0�����R�z��RA�O�B�h<�}���z0P�7#nU1w자���ĥ����8���J	"��b��jx8��< �;���E�yZ�
�E8{���{��`��ʡq�[�6"�`��7���z{W����Pc1z�J�x)������[��Jznΐ"�t�{��p� u�de-[�U
������(
2N�zv�Nuw
t����:�$_��/#Ĩ�$���u�?��e��y�0��ְ(���&F>��5!�'�Ҍ�P%y�"�� fr$�X���2%+�T�>�S�ݪ+�>�f0u�Cr��Ճr`��/Z�S��t�|Y���~Bb�IDo&��mTq��'�q�/���
r�ܤ6 �;��@!��Gd�:gt��Z����a��a��dF9�ܰ}���"�ۃ}��.r�3��.��֍��=>0O*���n;~W;Xxbs����o�T���)�`:dF[��D���1v�_E隤��^ڟ�Ί���<�I����
_7d��S�	c��1�à�+�RGK�O�/_�E���
qC�!q&'�c3e`��jQȼ˫�H�gǳ9m�#�Q�����a)�c��O>���$��V�W��O�{Y�d�9�4�)�E��P�Y�*3�n�)c�?:a@a�'}XPgff�3����*M�ި?��;r��D�#Ϊ�J�u~��N�8�,HX�9�O�
��|w��BG�r���
~�t'����?��[�kT���
��s��4����<�ణ���V��ZdԷВI,�r��)�R%P�
���R��9��\~/��Rs��=�c�ۄو�R�D�$�S����j�,eӷ]B��}�F��eK!�NL��P�Q�&��f�9�fBWǶM�>bs��VC � m����s��ӆ�F��7���c�d�lf�ɦ��]�j�3x%���1@6�:X\�?��2N
q},�������V�7>�B���{=%3Q��"�c���6��
�d�Ϟ\�R��(�'���)��x ������nxiJ�o??wF��>H�.>��WC�_�1D�y3�e�L!9g�6�ڬ���������m�uc⿂�C��Q�q����0(К;L��l��$�M�ͱ?�z@B��j��(_��u��K��K��Eb�5�f�0h�.D���v��;f�w��0�֝��H1��u���Oypat"��	��Ҫ����DYK+y
��[��e�1��㥌Z N�|+B1��]�I�_b;���;QHznu<1�,`r�����"K�JC���ʟ�D�����_�$ш壢O{ڣFFq����ט'��Q[*I�׌��s�xf��P�Hh�*>�,3�*�(;B(����_�;�OSX�LQ��ZT�݅>
s�����3C�+��S�8��`ǫc�}${\{��-�ů����&��L�7m���@�eXu�ebU|�QJTxV1V��������J�B'�Z�s��#e�y��c�c/�-O
�xq�g%�4<;���
�����R!�<.���*	�!;H�����-��!
��ڱ=zFs�@�Ŗ���l�`�`��C�s�z����G��+d�E\��oԯ�㮸�Ğ��=Rk�8eފ��^���g�*�Yyܬ�l��1�C�(a�ǚ�q�^3�u�����X�yy�+ǫ��+���p��Hq��&mV����o���13~��7���Q�-�<���4���@�#�8���R4�ҭp����H}v� ���|[^��L^����h�+�q֫���Ί�p��+'�c*_ٽ|�����}��z,����}�Z��٣Wx|�� k��<��WURD�ܵ����QN3z�4fE�)D-3��M�l�cᒝ�؛���J�S�fN7E�H7! �k��b��4Y$B�.�����Vp[G�<�'���,J�ʩu�v�^#'�ay�Ph5*J�̱R���-��	��Jv�ށP%�a�f�ŉB�%�]P�<�M��;L���6��dD�H��u~ވ\	��TѷR���w)t��=�X�Ȟ�<75&-��L�]f�ZЏ��Ζ]�]j,��Q=2�]�x�-}��߾��)U)@�_c��-O�v�Z�X�C�_zvE�K3�##Op�8�=��.�[��&����o�׉,��{rB�0g��-����-�:s
��E�ȇ�<�x���z�u!���M�Ԃh������T4�S )￴���}��xb�M���Z+a����V��cB]G��~�{�u��WZҾ�h����־���-�a��V��P���Wa.àlB��?�=�w�ӱ��߉Si�Pn�4鲈{� ^��^d9)�}_�qƳ$"\�L���_SN0�$��4+'P �����?�m�?���7+�&K#��[n_G�J��� a<Q�*OP`��8q�IK��{ ��Gzc�t��KN����JeG��	������5�����5�[ju���e�#��YO]��ڑ�M9�Ρ�����A��}_S��'�<<��]j��'��N�FA�� j�9�rۀa{V��ZY��r�kB��{��Ay [T�V����j%�^�5�o!���E���R�*��xUF�N�b�S{��Nu1�],�sz<Ey�0� ���_Te ���;��p�`߅d-!����^��\�t"rǈ�˒�CF�(�h�'#��V���|Ê�:#]�J��ޘO�[�*'���l~')p���H�k9�#�Xy|��CCԌ�H���+���Y���޶�}�yMj��9�q%^{F�f!0!�Tc$+�=��g��B"@!嶽w2~�̮���ߋ��+�@���샲�3U���Y�M��4A-U-�o��M��D�V�-��p��:ۜ!�Ev�}�;3�c>�]�ˈ�V?���K���-�X�0������m��N-�݉�(��)�b��w������k�Qe�����0nݴ �>�b��$�%Dqm��T<���<���=nL9DT$��A��vTwrJfF>�	i�>]�
I	c͕�j�������E��+Mަ��+š
��0a��'��H���k��������b/�1�8�6�[��^UdPYy��s?��Q���k��
�
:���X����t�{�?��v�g�'������d�N���)g�ś�(�r�˽q|J�3@��	���J��ϓ�cG_��R��V��~Bљ^n�Y�驃on���PE�ڭk���kAH�p���@S�N�I{���F£�mީ��˯�$�a����V7o��"��k�o�u�1�'��
���;�O>9!��mk�F0NC#�e��	;�@�\X&�ӑC)�]����_l��؆�զ�Q�3}�����/X�����Qx��Ȝ/�@l	��G�h��X�iԗ���M���j��t�Ct�\#�%�hN�)(�pks��s|��È@����Rk��#m�;GT���b��TvK%�m�_�Rԟ�"�{9y�P�%Y�^4�$x�vb:"���T�4$^�}D3���׈��1o"�g�,����bN���u��~�6W�<�='�d���to���g��
@XRA�w�=��}��M�!��E��<
|S�D�A�Ƨz�*>y��J^��M���w�mx�x0őÙ��J�=���_/�ϫ튯� �/��+��u�_A�$��#ߌ�1�q��rɐ=iu�0L:7�f�E��MAi;P�iV�G۟"ԓv�犆�ƭhi��d����;<������@a�./;�V���* ��?��HS�`Iw�R����*�dB|I�U/�^�J�7�E��/�l�aNJ�>�I-,�RU��-	̇1�\bp����?�S�9i��nn���O�)z��o)�}_�����ɹ�XR8j�\V�n[g�$�p	�ѝY	��ER5v3�?�P�vG�"��a˵�r)�H��e�N^�\c0俶]]�� ��$`�To�����~�7��8QX�G ��f�N��:��ʉ���A	��=4VJ��y6
��ݭ=/�N�*��)ٍ����N�\�ơ~�A����!�ku����3����j�����pb�~���.�w+_Rs��~���;4pS������u(}g��oRψtϊ@ڦKEr��(�wH�r���'j�k>g�3�a���E\���$�U�]��	���i�������Ck��m0����ش!>�����?V�f�:?hy�K�l[����>v)�S�/r����6���X��4��t �(j�6���w<�x�+zk��!�T��K���%���ġw��r�%�T������#/��.ZiШ���Iֆ5x˨?y�J��2��ML�z�,�E��E��%1hE�lU2�싿m��^B�BՔ��.-E:�eY�)�~{$�C��LB�{kn�&r�}�Lq0Γ�� 6�4�>�N�-��5���=�/#�Rf��f5ӣ�8K���Ē�Ԯ4�T՜��~�f�:i/��/笉�@��0�t��PFm>A�������0#f�"��97��v�8Py5$���#����W}\�)8A��I��4'8ͣ��1W�1<�#<��W `��k�p��زx���$A���!�y�������E;�|�򇛞�ʘV��X���o�L��Q�.r˞��(8�����2�Av���]����u���w|�-i�Z�*�HJS??B1�+�~�ْ.��u6B�9���e�p��M�H�8�^ײ�ˠ#QR&�QT� 2�.C��	�)���_X'���ؙ-��	�2tc�b�Iysp�����[$�� ~��=�~g_��s�::�_���jJ����+=:�k�J���L�U��l s.���E>��J���	�س��]��*S���<��V�'�/��[Q��`\83̌�%�j=��!���%���F_�V������p,��8_`b�<DÙx�[q̬<,,�eՍ�+�A�o�:�c�E�S�>���"h��c"�W\��W�g�y����_͉�!N���i28r`����;?�V@r�]6$�)���K;�����܀�6ܾ��G�
KK������8ת�����?���Z(�>}S�:�U���0���W�M9�����N����<�/��6K�]y�?P��2/ƨ�I�>I� �>�Iǥ1W���M��I�	e��O\��`�z#�h��wdZi���fV�O�\O�e��O��N-�v�&f�w@!���H�A���������wq��FW��V����V����&h�PMk0��+Nw����=9�UN��e�%�^��<����,�w9��ը��t��)X�j9����6ge����Q��"D�"��*I�RάV��ݺ��>�O��J"ʁ���X2,�p~�[o���{`�)}L��#�-�t���4�XCz��>i�aTc2�$���K��]�~v�>��c�!-�n��!�+�{���G�Rn�6�:�4
hy�˰��\l:��L&ή��e�E��`��~ H KE/�u3����K��V�������ݑ�2���i�ѽ�{Tx���w$�&�0�Y�$�9Jq0��Y[�K`�bID4N8؆N������8��~�)(W�ǡ7��ȃmj�d���Ou�3Z����HA�&I��禼C�O������IMq��j��"��n6A�CZ��m��a�;~SG��ja.3�3lE��-z�d�����I�)���/܇/�,�5�{�
{ŉ����դ�P�TU.�H�Z����Wiz���h��	�`dW�<��k���i~�6��ǐ�uJb��1� ���| U�
] ������֫�ʮc��i��ΐ���I�1�z�ŘA<�{�=%qA��tb7������×3c2�G����I7Û��G��r<A>������I�#ѵI���o�� K��� Y���y�� �cΘ��S ����q�Q�EE�0��T2�{���GV�'`Y�otS^��\r�ȝn4�*�Kȃ��gM�@��٠��qh.��m�fh�� �U�8j5T�S����!�kn|��[�NCE]	栁G�/��� �Au��|���6�b��4�y�]h.����z�*��ڟ��M�
H-8Ѿؖ����@��'���z3uy� k. ��6���5ݝ�!�o?	��LN,��"Zw{ؐӤ@�+���)��A|�C�������F�z�#���l)�J�$�k��
�|0�~�|p	ǵ� �|�����־>:�P���?&�^"AZ�*�}C��|�q)?x� �n.n��a{���g�<m�g	���Ý
xY���U]��r)��];�Q�M~���̬�����
��9GV�lH�6e0�(������1:���Cr2�Đ��LeC!����h"+a��� xeE��ޢ��.��Ί<3X&S�a"X��tI�b�L!�����X~�ml߇�G��J��kt�/�W��5V�*̲SҶA��P�J���t��C��Y*:{��Db����j�C�kk�U}ڦ<��6}z���sY�q	�򆆜T�	���B���M|9�v+����ڢ]���RMB���>���bY�Z|a�@��rަ�J�-9!d�	c�x���a�<=��Y/��=o���YO#�?�	d���>�V�ָvC��������4����Ȍwr�`C���TIBf��w(�+.����s��j��y�WT�6DQ�~n�i*D�|������tRY% �˛�3�k����@�=��%���l�.FM��#�����\%U�z0WH��m,���,A6��O1|p[����m6����6$Ģ�^����~J���l�+q���oa[�b�1Q)I*0!%cZ��X.ߜ1��k��ߺ�#"3�j�����41������+�GK�艶q�����j��ix�I���۸�m�!�[0:��.	ϟ�t�� ��3ɶNFc���V��/�8X�N����>i �"m�����ݹ��Ĕ�Wn�1� �K��D�r�����J%�`5���	YD�1��y��8;[	�V�Ye�_��Ro��ǩ����]Vij��>]�l������C����8��Ri�][�`}2�D���.u��x�����!���06����@��F"\��}P�M�2,��5Ξv��v��aT<R�s��(!o�W�����f7%;Ƽ^.�^��D�OHv��ar��Z���n#����xQ�BP�t �����	S�C�N?tY�1�^Ϸ)B]P3]Ϣ-km�R�kN�-��(R�q�p�<o	��>�����ø��#FS�Xl��p�؟yT~�6��������UgSW�����Z���[x�9eé��&�x�d���	=P�����djCU�ER%0!�]��~��e�]����Iߍ1��y�����D�>�	q��>�~�����Z�~�nKmK�g����iv_�
T[��ަ�ƔH�ϧ���J�.HZ�F4f�\7_��?�� |�pC�n�C&����)�9���q�̤�P�8��L|T�61k��׋�iB���w��
Jo�N|��k55)'K}�&�Em�]T(.�'�cf�� �4������ݡT��oMJ��ٸ*S��n�*���h1�[��dP���F�g�9��w�W��=���z@�>�]$���ļC���0�"q��h~*��bӛ�,9�5����c��k�^,���#�f��'ĴY�YE-HC����"?�a`yy½����,�TR�M8jHd7���g�eg�g�����ȩ���sC�g�>;�%�ը�Ga!^G��u[�	��J�P8���
R����VB,�-@f�����ŦG�b�x�d�9[�����OG�A�_�Ŧ&�L!�^��HON-a$�3p$�;�vIlw��h���>?Q�,���%�H�uj,�]��;ju5$��z����9I�l/��P�d�G]��g�'�6�3IV�$�-Ѻ�0�MF� 8�g8�������.��&HcL^UKheMh�3��H|l<7�#�͊�ݤ@+U�~f�-�����r`
�>m��5u�>?k��j~C�u.�~�0(�BS�d[ �N�O��s��%|�Y�F�S��Cc�/�X�,� �]�p$�Xz�d$Mz��_���� (��u����Q��KC%������Ξ��
���4`�����aT�Ra�}�V������d<�*-4�,H�Ё*����f��vʓ�9v����^����Չ"�q��0�{�6jxЧ��h~��%�R}�șa_�h� ���M^\� �-��D�a��4YQ<��@�f���?<��SĴ�7������0_�E��B$���u6��0n�o��efo
H�:O���n\L\d[}j�eH�2g
�`���+
�}VX8n��;��~x�u�-^(-�A���1+j���@ʧ⎋Xm"���ԕ^�vbν�N�Vs����$NQ��Y>Vd���~G���6;�^�cR��#"�p	�y�����#l,:����7�
��V+�B�ހ�P�iHpu�Y9�d��ɟf�:����]I�6�2L),���I ����+d=婱�`5tRjJnA/�MK� x�j3�Law�EL�ܩޞ�8����h[����K�Ni�>M�^:S"�!�4��7̭PKɀ�s��R0����C�b�uR>ɀҼ9ҝ
��k�ULgou��f�������8Q�ť6�u`���d��nHo���b�@ �z��K�v���R�@G��i����ߝ�g<�u(�>��5���9ǂ#迾�Un��z�S.��"r5��h{!e�GpϜ,!i�T����o��Z��,M������wj2�G�Ϭե���&�歸��]bN���]s��[�n7��ջ�dԓT5����'��V�@�W����`��BGV$�oSVD�	�:8����l[�~v2t���TAf\6�.?����Fe�b'��>��kˤ�
sW�y2���F�Q�����S���vN��<k�&gu=��Gw��ى8P��U)�-T+�T����\�}����`��Ӈ0o9"�LF�yգ�"����uNEJ�CRL�փz�~�S)�y`���Cڣ�ܳgB�\��<�~cv��P|E{y�&]�ߜx.�^9���	DS�aX�15�)6���$�(,��FT��!O����d�[�mb�XMi���!�(�J�S�&-�>��)�I�}�?���;���}ϡ-�ć�d�a߃9J��`i֏�|�{�5'������E��(|�� 3��f�9胬Z'ɶ,a=����pH���G�G���a��,�H���(Qժg1��6���N����3�-�3�0�=�#"�t���by��6D���t��Dv=$�W%��w7���G h-��L���Ir���D�&RQ�1��V`X�EB6C�C9�b�/h}�EjEG�e�.j��&��s%�E����{�$��.������/���vv��cN����~~�H�H{��A���v�.��]a�S�ٛrɠ�(��Ň��R[O$�t}���F5����`�%��Au����~�e,���Bk]�`������������ME"S3�#S33���BeH4��P��/jO������0�X��ܸ��8C:˺ u�A�y�q�4���e��GL�%;�X�˦�Mg9�sE�� ��0ݶ�_�-Ҕ�N)��/�1�qƓ"���gI�����#��M:<>����6m��{���=a�`���yl�@�Eˬ���'��u�F��4p����Cq|v����ɟ��.�eA..!�*|=�\'�a���� !�>���cK��C����;f�^�w.8#O�ܤ�ص����3���vϰJ$�Lw �ԣ/ly������Nv;u�23��P��
j�3'Q^�z���k���nN���}���X[��'�ru�N�9���Y�h.�ǜKS���ah�����T��H����O.O̶���N?�ӁEa4�'4}�n��t��{1���1*���|����8޼��;�h� ��CsՐ��]����Vi�W_g�4�*��ۓ� Gȳ���~sd�P3L(}���j����EQa��7Y���tޫ�ar0;r)����ō;�o���?2(=�[(��KM}e�C����;c��TS��v�[N:(��v6Ŀ�Q��&�c�g+6Q��u�a���F��ԭ�������3��M��>�h���m����iyY�F�?�	^���	�	�f����9��WC��zXh�W�I�^�t��8"�9�]Կ�-Qr�u�V�Ą��A䟯�wjm�?\ȳ�x[�iP��1�AM[��(��43��4Y�(��K���&MVӮ���k#AȞ���ex�2 ��E .�4��Q3KXW�K���c����D\�\�^>!�� ��<p���O����B_�diˎ�0�����FT7)��(�k�pd	~H��o��D
�����e��;� Q��b�rgA+5 �.��9i������PxҒ�Oq"����N�*���FA��Z}�t���w[��Aa.�u�_��{sS�z{�v7=��Ϣ�7J	�uX�!8_��iY�N���H(&�g�
���X���0Ƶ�Bӆp���N�go���pnA���<jL �s��?���u}�<��ۿ�P�j�L5�8�z�+~ʾW��14�$���5S�5��W���#��Ⱦ�ɉ��&�Od&�ض�0�>5KQ�O�/������o�:���g\l�=q��3<t�̋����h9�ɨ jx��"[RI�q-�_���Oe-�
Z;����x[�uN�A��o��6�����k��k�_�`���Q-�!A�Ӓ��ZvACW�!�pv�C�D'F�~�	�ف�Iz
�X����@���׻�M�8�
�K"4��E����}wT�� Ȑ>����G�h��Lh�\��"�ag��ҤxF�Z��
��B��+R��'p=KΫ���*8���:1PJv2�+�eG����צy���vl�O*JBR���t�O%�t�ʴE���t�a�Цf R,x�%����.B���u?Yf��G8�^Řǰ)��!{9CW�dngS�����@�#����8w�ɕ<��I�����ne4v���,8C��=���[�i���G"P�	�I�5�5Y9��&`Jg p������wV(<�k�]�+{�*8)�F	�!&��L�p������)��rZW�W��q�BK�p6sE5j,:����#����c�B����m�� ����7�K�↠_+�g�jn���	�P��M�檈�!�D.�.���-�\W`�eN�=*���QQP�?���C���mi��,�
~}!��A�_9(���hư�v����1)�A&�TP�����=!���pb#^����|��C'�vv�A�f����r
�e�(G�� �0���I6�V�ey �1f-� ����f�@�킓�����G�lestIB�Oִ�|X�n��zH�K���!6�i�Uw5���6�ݬQ����{/�4B�V�}�X��x�[��n����kFW�%�����&z$h �h�aɳ`�?ȒImNxr�9) ����ጞ�2X���F�ʀ{���Y���O퐵Tg�]԰+��p�NJ/��;��	�d��
�uQ����J���,� �+�J���~~��Z�荬T�P��W�*����Y�p���$��dy����Dޙ/�1�)s���zN�-r��re�y^o�͡��f��[n��Ϭ��*����,�8�@�E35-�d�m$D��n���Y�������0Z�-�N�H�Л�\�t�h� |�*L��#�ˍR]��h��^P�e�E(�-c[�����͒�GP����	P�FW�3��c/�f¤��p�.PT��[�����"�z�9��� \�MӈS���R�[i)zV��d~
���2$=�
vF�Nt�W�!����4�Ig]��5��w��m?��g��&�/�@��7�9�S|�_[�	�w�N�P{J��D93���Z�"��M����מ?2�vF�4�7dV�(���Û�={��S��4�MK��]ֶᾙ`ˡ&��y�(���S� ؒW���tF���P�����SG��KR���#��|C+:�O����kt��~�=���؄��	���f��p�3��l��i'���et�FkI�S�P���d�	�_����D��]l�a�ְ�+��G�$��B��.\o$��{�ܗ�Y��U����)�0�����&��,Mg䶨ڋ�Eb��?��WN�q���L93@����U!H���#�����Mk'!$|�p��j�w��6<�t'�#�	���f��r2b�A�"dS���B�������l�S�XS.|7�]~��ٛ�EVGʍ烔b��׹U�-��4| p�Q�ѹ>( '��$5#-{�n5�c��|7b̢�i�s�*�L�������4Z�e{���+i��>�L��׎+����OBju�		/�:A�;���U���ǖ9��-ǫ�B�7l����B��CV�س"��U�)���H�3�	�Ӿ���㑛�y�i�M�3f@yU�=�˱�Tƥ�	�I��%��P{�(��"�`)sg� g	'�q��|�� �Y)N:}��QJ:��N�u{�V�f���}ۍ��V���r�h�!N�uw�+ T��Y��Xa�d��4a�:�ڀ�1z1�
��:�
�>��:J��z<TŽ�շ�Y�٭�HA9˚
�֑S���R��!��ErC�>^��x���q��9j��kWt'��Sv��
k8xJi��cBB#+�~�m�� ���K��׹|P�̈́�3ulږ���iN59���tm���7�q�4���!�O1��|�QExy5�uަF��66Ȼ���<�+C����2p�����@/�$���Fx����0�S(d�jH�Xg�X2���2gy��5�c�ȸ��uX����YdC��V�ȕ{��u�TI�d�YR�m��EZt��_�����(�LH�~/!?8�� �sI�������g' < v��7RR�p˝���c�Ɛf�\��F�8:}O���
��L���*��r�L�������q���ߪT���Z��=FI�ߐw:v���j� ���n(���b�����*���iZ�&zpv�Tc�"~.�`jr��j��ؙ#:�o���ϝ������4A<�d�MU#�Gv#�m�h��nޯR[z�	�ǐ�@G����Xa� k�Y�&�6�o
��_��.�F�pdcq�q�B�ux
�/	���)5��hF��		�ҾC��򓅎��C���D����L(_i�>������V��%���տ|.�`�5���l��6e���s�~@����~1k;W� �%y��
���D(U���U���5O��XA�Vf�����Am�|���do�$���6��M��>����n"���Ac2e��"��Q?�]n$�]9#([�uRj9�$
�қ[)wk �3�p�sbD#!�v��3�0m���6�z��gK{�F���}\��w*AP�3�L����a�Qq���(1u�B�%kQ�C��ZgG��uY��M�S�*j�m�}����7��C���h][7��p:7kg�-R�X�,C��-b��;�4Ny]�sG�ۈ���K.!z��;1?�diX��<�l�/��π���5���.S��h�>�{-� �f��t�ߧ�䅘����/�����3ӻ��mmXNx)�F[��b�>:��Ҫ8!hjXP67�IF��u/�u��^rf����}��u����\�˦zpB��i}h��mF�w���a�^e�D�jp2�3jt�
mFQ/��@�6#�9>��#�"�1C�����G���;�^c��~f~Ρt����2���BJ|d��M":� ��O����l ɸ��s��I�}%�Z�������m@��<��T� �[����<$]cwX�P�_[G##�ĉ�Nμ@u3�%�1EZSJ�ʺ��}d/s>�؂�M������j	�#��?�����ƿ���A�	r��zUJ���s ۿ�C��05�����r�V3�������aQZ�-8.�R��S� ֖�buX��i*�2#<u}{����8Q�`�
9=&��4G8��*�r
��[�N�h�� � O'�x�'�|���;KÇY����d��^��~����$�iFf�orc}� JL���N�B{��gwX�x�˓�:�\p���n��)�$ғ�{]�p!N�k���7Ц]si��cK�;�FުQ7�G��=��3���2й�ϒ����I�ud����]y�n-�B����ruT��\dj,3�Iy�b����K�������6��|��ι�pRk���}���^�\e��gY��m3{p�L-*�E��l~�R��� {��^��?v8Q0Z����a���ǜ��Y��$BJ��i6�t�X��^����ʹ�e�6NՀ��&ø[�x��}��s�ͬ Y#��Ti�� ��P5�Imȵ�pK:3���G���ߚ�	�,����H	>_�=���Fɏ\^!�j%V��i�����p�,~����õ���3�U@y\�8�M��ql|`���(�Q�:���:�z�|,����w@�cN��N#���څ���cQȱ�^nz�/5r��6�z���6��o�5O�j��z�i+��GY����?���D��].D�}`8�K�2�bf�Vb�������>�1ЂW�RF��tp�OԄYC����/�׈o���t�6�ȋ� Q�ᔯm�k���몘D
ٟ�o����D҃��L�[b����zu�B���\����=�\n[��w������W�bT�d3��˝0�Qo��zm��	��
�*�~��x��7�*i�������1��Y���u:</��񒄧��5젧 =�N�-�w}eD$�ܚZ����H��C���B{���48?zy	 �|�m.�N9f	 ��)�9?�5���ek�a����
¸1H  g��fQ4��Z=����M2�hY�yؐK���
�:�>?��[���@SC���t8���!�l8����c~�Tד}k| ��­xY~�ؐh�*_Dh̿H��c�u��6�´�%;��.[TxR�QK�iH%�E�Nl����G.\���O\�I��u=k�o���AF{��y�2##8���.�aU��s�ɣ���eou����L%|	���%�r�j#�j�u>�yŬ)� �km�~�o.R��y�T�32�ϝ�'JS��Q���ȼ���Պ�Xl�Gn�,�L�D��4{�1*������_��[�å�{�Eë@ 
T(�^Om�W��<����_��5Q�G\�������x�N;�
"�o�k�������ɡ���j-���$9)د�G���/��D��lu�v�IU/��B�=����ET��;}
�B1��x��@d�&�6�,�@=��P�d��j_��D��2����WWJ�f���
�5=)���#�����ۼ
�{�]�t�x<X�$J�Tl��,�����>��0��	`#L/s�߼^��Э�G���| YN�0b�� �q�Vc�l�*�$���ؽ�`"&���[�r��j�p�"�?�~���M��j���Vk���S pj;�� /a�S|�Y#�δt��� ��`���%0u�=�_q��
�Mu�?�&�g��}���7��D���h��g�^A�0�pn��(��-ao��vk� d��ٶ���N�t$ߓ9K�og!W����=�<�����?��>%6��x�w ����L�a����#�!Q��V�5�3�w�r�:j9lLhQ��8J���1Š?:����N��M���O���dc� �|� ���)!Q1�,�g;���.�r��Y�85j��ߠ�ѳ>����8���>���=L���ྍ�����,(x�f.hƭ Ʋ؂�i�M
�P6nߥ�ڶ��(���8ftgR�c�4�=JD����o�*���F��)F���2 ��6��2�X���{�0Ě��yS��I˶u�J�:���?S���*p��j�z���]�e� �B�?�?��"���9�)���
�L�/�K�*\+�FC�������� ,S�kl$�%�)}����Jz'��N�g���������S s�K�ޭ`��.̔0#_W��7��1�rw�i�zCc�C&�`�R���Bu����x��k���>��L3}���"�C|�h�[ΨUv J���`
Rj��3�j\ �L�^t:���c�����ߺ���Q��ʎ	��W��*�<Z�$QU��Y��u?�U����[u�DǋT$*�\z��{��l��M̤(�:��;�4