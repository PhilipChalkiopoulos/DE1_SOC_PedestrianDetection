��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z��4֬��9�A��;Un��Gh[�����<�#�L�-8�o����X0v�c�4��S�`U��� ik�{=�g]�C�+a
>kN}%]q�]���g��k���Y1��Ǟ�H� �a�C��O�m��� ���:G��ᵑqZ��6��i��[0*א���H��5�|^DB��xc����>���♍�@�Vq���2@/��U�_�6ӴsV|���h�ßXCp�s�����?�׾��Y�0�č8�y��V;���ϥ(�ֺX!pR]�n�Y�#m�IR��C�[Ѵ�hӽ�ޞ�8�O�$�7��s��dk{)�Y��*��x��\�itRFD�~�2���6}
G2q6��}�qJ{��|��T8qlX�8m���6�����rRmP���愅�ʦ�_�~�������,�aS�Hv8Y���<I�%�����$(��|�M�̗�T�i��'rYciˠ�� �Xn�Z�������޸� �ï�SO��g�N�d(B��}G��|Fr����RMJ =����c��ۊ ��PIw�DF�o:P�t���N̬��Yt0��#��d�� �v"8'�0V�ǋH~� �,�P7�9b�zb�&ӄ���7l�3�V��{wC�=� :T���4��Lq�TȀ����"�vy�Ri3��g`_]��H�C�)���bli�{�40?�l��s����b4�t}�������b�	a�);���T��V�p�����O9���<�M�_��1n�+���Z��0p��v���#��u���_����cE"��{����3oL��� -�N��ά#u~j��J��F�i��Y����03����-ǿQ��^���G�����Z�;^pi6Yw� =���e��Ď.�s\�.�`}5�O�:������3[Oج���N��?�!����mf��.ö��lss5 ��x�Ҕw�g�XxS�/Z>�>��z���s��u�.�-۾�7S�x{I��Q?I�1�������`':C����_��;e ��w"=e�=y��&�����c%�13�.'޺+���@���_zO����:zAC�"L�]Cx$u���!jT���\b�v�-!�#����
�r�e�bܾS�ҁ'��!ѵ8@�X�A�9�!�}D�nhW8=�!����Zx% ��_\ϒ#�]��ts�!(�ӧ�Tf��A��H��uN��)u	��]�,F3� 9q�J��ƩX4�f`�F����(�;F[�>�/�q�Ʋ��9��ܲv���I1�v�㜏_wԱ.r��o�E�(B���YJ�J;\�B>�m����`��e2�����^�y�3>��9l��7W�Ç�Q�����0mǸnk�A��u��py�?���O�mC�_�y��oX�TY��um�V�����Q:�"��j���D��ƕZ�D��p��V�54�k5�f}��M��5�ˤ���<���y��o	$�}�XFP�%K~� 4������26z���G����Rh�b� �|�<��*�K�֪�(�k��R ����;�̦�C�>G2���Û�ܔC�C���XMW6S�ʭ��lh6�Hbk�8M�2� Pg��̾T�NӉh��YrS���\_ E�g�����a{2Ȃ����TMNU�-��4���)
=NWh�3\����4R�7�C�a�ށ�BD(����m���
=^W�P�ݤ�|P�2�:/�S0�䙴��s��r�7:�0k�f����^�&t��,70���$+Q�\.�o%�M�	wؐ�"��ǳ~��q�G[�XIz!A����Gj���^�t[��S	w��m�AB���kL�!(Ab�c��K����xh�AR�m�)���୧X�X�b���OR@m�3[���էϠ���� Z����ذIQ
�pX]���XR�
",Up���m�m�3�#���E���o�s���M�Q���à,��{˴`�݅�������E���@��xi���;���߆3k{���Gx���E��xH=�����EV.�d}g��lU�Mj���Oɺ�_%1P�c��m���cϓ0��;U}���-'E`7Q�?<󊈁JG�'պ[���l}#)$����'B�B�J:�MH�l��HS9�{�t������7�L���^!��XE&4/��IϪ��!h�~�↳S%��M,����E��L��63n�R��S�϶�S�*ëM����=��>��}��k\Q>Ըg:0�%��y;�8�����CAdmI�5����%��Ǫ��?���]l
����8T��R��p"��*M����/�YX
����C�3������
=4:OX;�.�t�K|�h��8�Êiy���5p���`���:��J��9�rS*�wd�' ${�)p�-�i�A�'�^�@�"��yub��}����kx��,1�f�b4�ɀh=�; J�P�ω�`�����PF�ȹ��n�$Ƣ��X��u��5;�gF"X�*���gg�fJ���8�?R�@�3{�qxs�z#�R�68�(MC2O�4��B-yJ���	�Vr��nL4^��r4�|�M�[״����:c�f1ŊvҩH3!|�ӎ��0�,�`Yx�Rs�7�H�lI�W�A-��ˢݝ�d� ��:ȍR<�:V�����6�� �&����w�����L\��FD��8�(z%�U�P��"��<�'X��~�J�T��hWP�
+��(FV$�'�G�n|��UsR�p����)�[���� �F�q�2��ϧ�݅.g�߹�ˈ
������׳ ނX�]s�{�������o~��z�ŉPV� �tM�GG�?�(L� �|A8�^��*T��ϴ��Ջ��`�4�P���G4�=��`�:W�����
�U
0^ۓ�S�/2���	���>R;��Q*t8�A�&YBd�r��������� �hj�� ��R�m�Zj�r�t����SQ1��6Ҽb��h�/(|�+�5
�F�]�J}̇6v��/P���'u�|��1|ސ���ơ<uq�2�-�K\�\km U�ږ�w����f�(�q&��Ds%�<d�}A�o����rq�̀���A�H�f�����Kv�)j�fsd����(�<����!�AW�G����cxQ��:>��<��z D&]������i'<�w�}�i6ƙ4�\���<L�>��I�_�P���Q���_N3͈1H̻���m�K*CƩ��� ��8��t��?��X�x�|�[����H~ ��NP_�֯aS�M���Q1����ܔ���ϲ�7*�x��oPM.�c���~�f�/���9<i�9������}>:'5q��q����!�f$�E��r��h�s�	����'~Xj�5;Ε�Yˀ����� ��Z�L%�S���2�`Lq
k��-�]������]�=~T��ؤ7VΕV�~?��GUڄc��[��$7�AJ�e'�äU[\���` �>�b)��K���Q�c��6rve��EJ�;��f���&mK@��;������3J-�/���^�uM�8��H��w��Y�;`B�Ǚ%�ys���YO����s8`���	�U'X��$����ɍ3�/4;[E�������/P�$=��{��n}l��U���v>k�Ħs� �df/��\3S���;v�������*!ָg��0���t>���������7�����*m��}a���Y��T�*�=�c��4�k�,�#�c�y��ϼL��lgL��x��D��}j��x�n�*��w�S�PDMȰk)hX:�Ԡ�i����o��w�(a�&o��� � *��6��1&����&��@*�����s�"Tަz�f��|SkQ:���%� �jG��L�0��+o�O(u���$�2#D��K���}>!C���E��V�ƏΡ=|�"�a>zR�	���������MoW<�=HD����bl;~8#(R-��₵>,w���c��.w)C��4��2h��>�(��������R�8:ݹ�bx�?V�,@�\��>���<GK�Xd�넡y;�o�$��=�?꼇��E�=�>��5l��]�І��%0%X�h`bX��+]ČRWV'���.�S�O�������\ԯ���RA�O%��}�����g�<ۚj}��O��(�'���uv�뇋�-����~��/l����+�6�+�X�!��`p���e�4�j��՛U�as^�<�7{_�m�HZ�`�!�C��b^�&w�ǥv:��Y��<m�*� ��vn�I���bZP��X��}}B4=��Mcu��#��<��T��&�6W+��$�.����>��Y��b�J^)����/o%��WA�
a�<��3+�/\��^!�����mE�%%c�S�%|�9C�Y|�T�O&�A	e�G�S]�3�����Ԟ�F�b��`":�5:���<�S^jl�Vz"��B��jSȕ��rt�5���9J�IR� 2V��?�s1�"�}�m$	�y�\��� ��n,w
�OV��{�G4��f��Rȶ1�۲AQݿe q�v�,��~g�3><���.m{G�����`%�]Y���������~[o����[��Y��=�S&�E��o;uEQ��gnD`�n)����qI������Z�j�}ަ�\��8H셤 ��dZ?j)t�U���0�Q`�RS��������LPxq��$)�a��x���x[�T>ʹ��&x,V����M�K^YI�>�.��q`��KZKĀ9���hIY�,��׽���R��y9+xh��ro��	�O�u0�c�nnF���T��cz@5��h���,� 40���7w�xI�}ao�rK~n�`�u�ǉ�?������GG�L����.��jP��t���!���sl2ʺ���OY�7z��1��3�ބ[�����=V@��v���΅����|bq ��@H�o1/��J ��*D�HwÖ��͏������bw!��|�뗚jR,@\�F����C��tk�N�AѶcP"+u�����Y=�Ҍ�������*@��aQ
���F��]F��~�e�қe�� �"�������?S;��f��ϸۆa<��sg�H��<'<�T	A�J%�\L�{����k �o#1S�ڻ���������C�������rُC���u#:��{Kc�(�r�y��[�_�m��l��\8U嫛c��g�[ '�<�oy_H��"bS���%��A�\���c�%J��?Y��	 �;��-S��C ��w�z;�6��H.��Ź�R�E�I#{�VT{�<��`P�b`!�~�� �F��-�Z�D��-h��Gt��i��N�A�>Xj�R����N���aE(k��z_�7*ʁ�÷_}�U\y�g}���''�&�d���\��Y���hI+������� �j���	�K��:��\�%�շD�a��1FmjB`D:���z�[
(�Bn�\���=��wQIap6?���j�54.Epw`g�!Z��w�!�4a0W��'r)Qe'�6�y.������FkS�xk����
��C3���-3�*ifZ�8$ G5��H�
�3My�	����Ֆ���Z�KնJ� ���l��|���}�j�c��h�!\Ze���D��V�B�\�^(l��Ԩ�f�����8��nEA!Sޝ��q��'e��7ڹ.e3�G���H|_A����o�V>���딩�P���4����(mv���X26[7C����eO
���d.�=��6Ӫy�k���
ɵA^�m)�V1��OBO ̯�R��Q�B�~���'m�Tr�q���h~�O5�x�>�h�Btt�Q����G�Y�����sh^���B�?�����D��w4�G|
S>� +yB�8�B�eG��g�e�A�� ��Bg3` ����i��I�<�F��M�$�ܯ�ɑ]6ҡ!"n$wP��*msh��)c8?"�lu{d����˽0*�-N�v<m:��:N�1�������1��$�N��'�u��%�)KY׬�<)�S��v��Ac;��������'���Ld_&?��J��pW]���o��	C��b����J���,�A���Kf�꿙��(W��J�*l}�Y�#��͆}�~^NƇ�}0�r��؊QM�.�J�z��}�x%~����{,�A�`�����[f�[h��Cφ:�F�Ą-3�/���+-$ڃ�i%@��w8����!8�#gj�,Xb֤h���5���%E0i��K5������K�Π��Cph"�&�M��Ͳfӕ?�)�0[�����>�� ���ΦI�3h�)_�����.������֩|s�*��5	��v�v���Sn�(�DL��ϯ��Mga���'���f����|�B��+�X��GMR2����#�h�D�Ĩ�_�r:4̕��R�a�8��;&�(�W�{�l|�y^ԯ92F�,���9 ��Js��"���k+��V�lG�ł�	�_|���]\�잻��4�:d��}Ȱ�ҊtH'�X���e�h����I�^Ҷ��>�rVߠi:RQ+�����r�[d_{��H�?�vQ���*��$���
���u����FE�0��JSslh����9��f��A�T=ԍ����c`<y0�˜�.��5����Q�0#�犏So�X��H�k;W��BooWL�+$�ۇ;�h����	��uook���RH@]�}��w�-�'��[��ۇI���XU}O;��S� �f��.>�5��3�4߆�.|��vH�=��H$�,����L})ʺ�yթ�=J����|��ЦR�a�ׅ�PvE��5/��Y��AH�v�2H �B5_3{r���暛q�ō�0G6b��<�|��<�xu8p���j�|��i���N���L/<t�黊����f�Ĳ0��u�+��6r�����l��U)���;b���=���UI+ny�����Mʌ����=��Ml�sF� �����_���}��f�)6���G�ca�l�$$�c�hr������+vcE�\�mT�,��<�+'��D�(�Ԉ|,$anG(p��F������f��8R�<�Q�W0�T�i�-Þ��R6;9(�����0�aИ�s�48|�6��\i�5�3�&5F��0m��9i1yb|0�A�F��Z�9��ƛ>�&�V8�T�9H�toO�ݐI���f���#cA.�������S�u����t��b�Ͻ����z��L�c]]�k��#�z�(AG�s��{��$ڽ�c�p�p���W�E�3}+M�E+��m���Λ�Y<�3�i�]��l*�t Ax>SSEY+�ko))��A��Ƿ�ˀ�&�Su�΍l2>�<�t>�%�i��ʽ���.�Z�#v��16A�G�1�x�,�W�eͅY�L�.)�I.��&���î]B2!���n=l��Tw��a 1��1²���o�M+�� ��ߡx�4���&�xta����7JvUE�a%2_Y`�y�Q�GD�l�����(!�2��j�ۗ��Wx�4�=�J�Y�~x��r��]�%[Ӿ�<�ڨW���Fv�����G�Cؔ<X��Qd2M)�~��O��i x��a�|��ō��:)��b�}��m�>Zߧ/�	�a��3N���z�)��	p��� ��Cf�A?��w	KgP�;U�/)>���D���;�9{�D;~��YǙBM��!�<�����#Hj~��/�;��G�Q��TZ�H����.oӏ	���Ĵ���C_������T^�!��u`�<��9ƬM�Q��2�~��~�Ǹ�k3���2i�b��f_�5���)���ӈz���ǜh��G��.,e�L�c�$D=Ym���G�h�Der���DR�=d���dPX�A��k�Po�Cm#�	��/��؄ZR�rR{�x�64����#ŐFr�&lRq�ۚ;�d�&�٠��3:#�3��L@�ރ<53k>������z��yu^j�e������>"��`��6eP~y�/<v���ۯ�(�Dĉ]-djr > �8� �\��?�3��訋[�� �\%��a�Z$���U�Z����j��7_e�m$QW) ���۟H�t��6.�iK�nS��� �MDb,Q�w�ұƐ����G���1ߢ�t�H:L�z��#��4ɼ;��az��b� U08�RY�@�b����-	K7-�/w�!l�
R�u�?7��䀤3ڝ�f�3G{��XL��y^\�t�V�_�5��*�ΨXm��E����߷ª���) I��70��7!?J���}6ںQR��zT	�tj�*��α�p�څ�V��ن�5�ݛ^����=�az���9�j�-���?���e$�9D�Nߴy���{f�>q)N�|<��5�F���<��Uy�f���Z[22�o!7HL�?�8�*#�b��Fq͑��m��MQЁ�n��w��a��Th�x]ȷ�>*?�@y���I����<��] CQ|&%�"��F0E�z��Ȣ��P%�2M� +�J�$PG���/������y�{�/sąB��,������Dm1Y��R�P��y�w(�����zL�v��z�wl�"_�^5D�a��f�o�u����}�/�j> ݾOեzjp	C�sg��������;�y[{�����J	���������+R`�<M~�L�~�-v4�/�T�CB�Avˌ��~�+��>VL�Dو�E�Ť,)X����"�Dv;�Ϗ�|�gSBT$�T�'x�o<�+҉H���~8�'ٝAxx��m3܎`�e9�F��4����>����H�i�y�Х��'�'�@��w��	O �-������J}yw����X||㽚������
QP_�rO�@�`.~CU��AO����tC���p\iݏ.@o���i\�Z�l���#���Ѵ�n~���۬-��<-mBU.b=6����i�~��V�Y��E�X~;�P�|_�?~]Qױc%ѩ.qS��@�sP�ꎿ �ϟ���P�?�����*A��2)=�����of�n(x�B�i�1�\�9A��r�?_��kO)y�����?�G#��-�%�OxMP�L=_�l�E�[����s{�8Z��t�Eo�_Gw�3�CC�%��23�<g�~�@SD�s}�F�=��#+�g;���"{jyF, �)�u�vu����&t��~�ȥ=ٌ� ��i�.k�nwэ=�;�x�7�!�,�U)��\��J|�u����䦵���G4��&=bt�x0�L��ىq[��j�84��#�Jh�N^�ق+&���Qf��5a�ߔ��M~i�z}J��7���������('��~/<�C:�܏߾K?�7|���4N��%�j+ê� e"���.&,�7�b�v����%�Ϙ���3�m	{��ᨃ�S�`Xv��"��	��$V�}�%��N�	�~F����1Iw�5D�K9���������8�
�n��l��%Elc�TclbU;X�/�����]�k�K��4���������Z!���h�ۢ����AaD�)5�ND�D���B�'F
5�b:�mI`���TҦ�>|RW�TǺ�>�h��%��߫_9�\qÁ���4Ӳ��m��Ro�/�Gώ"�ӕI��@2=�d-&����d���7��P��-{��q�\�RE�j����Q�Ak�$|	B�Y=��X��'��^�B�{hñua��ϣ�$���D�Ob��^�;Հ�Tp�֘ �������j�����d�sI_Ҙ(�h��k���V�Ck�#���;����(Օ��?��$�7H�oj�TH;�x����T�]�ۻX��'�6��{��X��ߝK������V<���#u��`Aɡ�gw�yW7�۞ibl�Qo�O}J�D �����Ɋ��yTwv)T�?,�2��y�ltr��$me���e�E�*E��%�D4���^�Kn*/R5:E����V��t����̌���_���!�	�M��*����DK�kڕv�S�<g�u �|�LY�2⽑�����	��Vf�Λ��Dɥ�����fM�a����<�!�����Ыo��Cz��ٶm�f+��y_;i`�����P�e�!��~v5=5J�jn�qCo�����#�_���	QqG'��F�#(2�Ҹ>4��	8��X�y�%vk8�+>im C�U�������p1��(�H@b��9��ڶ�`Q�A�P���e���f��a��	�R�p�HL9�(1Pk��hF���&���*���o�8��K9��u��JQ���^�2��;�jd*9Jӳ���ΧG�R��<x����g`oEv�P��a �:2�>�Uw9�o�5��.��s�l#K���|-�h�z���� �4q���q[��8���|lӝ>mu��EUU
P���2�������ΓYS�N7PQ�����j��t��y�8r��3'��<}���vl9�B{B&����D�B/��`����n���2�T���5`��t�|��:LT9W�g�ݥW&�ӕZ�?8x2;���$�hMo�6b��Έ����D[-Nb6���:����20l�����=�h�7���<䌍��ZM�롔�t
{���-��*s6�]�Eh�ިFb��p/�.� 0q�:nt�T5>E	�=���B��9���e�+���k�oq�X�y7`虶l*�N�s`�s�}1��r77U���㠽m�v��>�T��G3��O�=���{[¹Mg�F*����"�gD۬�[^i�4��(�-9�A���eZR��:���\_�@e��g�۸lNX��K�sậ��������&F�&|1��v�:���Z��N�����z���w��\��������Td0���xYq0�A_ЋP�m�7^���Ш@E��Ol�0�vg��951��OQ1�NCc����8K�XѶ������WLN�[�̬�c�~�ڬ���gAN�u.���"yԗV�
x�f�C�|<1�V�W�?��ރ�@��@ʓO6k���o�i����vUF����<�ѶV�!.[ih n'�c�FT�s�
h�1P�V��fq�o��[n&�6n/'L�Y"j�� ]��k��&��6W�Ρ���]��K�q�s�N�+Eq�]�^���;�}Yh(�^,��r��Mс�,A�hȏ�b���Q)��%壱U[|Z$�7�<�����ͳn��}�z]r�z��{^���9@�D�<j�yc:�����-��|��b��u�,��Q�\Q0F�+����/����RپI�o-Ӯ+�jAӽsN�f��iN�� ���9�����nR��U[7�D�,��gW��nZ�h��"�
A��eQ:������'by{A#�Kp�0:3ԋt���AK�*���@s�fY��=��p����//;=>��Π��l!e1]k�*-~p��a��
'�����ߖ��}aw��7R�WJ������f ]������ L@��J���'Z~�� <�B����<�6��/o�V`W���� ����C�ʾ�>�D��D��x��������'���{��T;��k� n����c��w�Q�MP��(��x(a�%u�0�>H�H�����;�7��BT:���TN�mP��2��Y3��:E8��E@'��Z�W���w\L���zx�
��*��]���ڄF,���:k�l"�F��X�'RZ.�/ʥv��$��׿x8�g؄�$�����|�U�/z��x#�����M�{���'N:���\�'Ң�M�b&
x4���1���8���V*��5�ȝe�zS�7cQǷ��!gO ��8�^���)���?�Yd��J�
��:�lp^ߊ�]0����i��a����L�>QXJ���b�ÿ���r"�����~N��^P�9U�O��T�B �Z^�����y7P�ӁU�
��/�� ���Å�}Ƅ�'VT��`�t��u���eg_�ͦD�)�3�V���䚁鿅a[Ҥ�|*t<�� ���Cj�O;�a��#h������bә����(h2��<ق�A�#u���q�iN�g��Cث�1g ^�1�Hyڛ�G9�pl'AԐڵ9��_�Լq�ge��Mj�%��+�l���`W5_����C$!D��NUe���rδ iZ��m��h-�ɇ��s@�zm"|Jl4=�a�ۙ�:���"i��z8c�]��RA*����|��%��/a��=h�Ԍ>j��^xwZ3�֞��.��̜��8�4;�TC#ШjCY
�[�<b�L�ƕpA��z���༾�#��ñJ�y|p�N� ��
[����c��B�X�&H_�Q�w+��/{��Sy�����?[���(N�mz��ߤ�GBx�M�3�m���9�
����8QL��Y��h�f�й�xO-���%��t���,��?:�A�I��������'D ����F�`<�P���qG+t{��,�Ʃ=H珗��I[�}�d�T "�w)�Q0XKg���Gz �m,�� �����o�s"?r�h��`��qfb��6���	ʔ�,���p����Ns�1�69]G{��3������	�E��G>�Kyoó���M��a��7�<kz30G2��MK=J"�}�k݋��R8_����$!�?��T���H�U+�e�����ϒ�1b	G�L^��E8X!m��'ܘԒ��実-6S�v8���Tov�LX�����v*6��`k(��CU^"�wV�1�2k�I�_�\Vdѐ�)��8�J�,����ٟNo��5��i�OD8����ć��p��0�#10.�J/Ҿ�p˱��?�o^�)�`�1�p �8�.H|Zp�p�֖������9Ϟ������Iʳ�Q�
_��)�\�I��g�S�F����I�?�SR2[��
�S)�c��r���3-�fa��H�0�@�P�[����FGc8�~񪙹��o��`��+ͷx�4n 7�S�� _��K'^*���Z��(�A'2d�7S�I0<��Q�H4����iT8>枸�������q�I[̌�����u�0��mϷ<��^���0�I���X�����ú~����fS��D�au܈�y�W|�`�zzF��WCs���o��i2D �;��ӿ�T�D{��n
�H�������8�j�S ٿ��7����M�)	4ܪ�;������T��i�;j�B��qDM��)XA܆
�$6�|�Q�
��b㪹�%�,��I]���x����IA'U��krY�}'���½3�9k�Ր��0�
D����x}Y!5יN����l����8ߙ���>$�+���D!���AA�n"�FN@�Oe韚���n�R��;s����GG+\�o0|��5�k�
���;��ʜ������U�5�\�f3 A/�Gk���&#NIh�	�C����UƮQ��,����=%���f�TV����M�5v")���*ёh��Ǌ'��Csr	�B��ڼ_�9q�tiEB��j0�l�I�g��3V ���ӭ>���	]q���������!�!�I�������S�����$�q�%�3���CM�yO�,:�����V�ծ�4�07�<��^9Sj��u'�N���ђ�t��L7�î�B��Y�~���K�,�{u�#L������oԸ^�2A�s�V���k���B�3I{�3)�1�����#���E�ߟ�M�ub��2��8��/�]u���p`:ְH�F�'��jޱ\�(27Ŵ�8$��㱓@HUxe>�ٵ�d��ad{_9�fC��$2�ϵ�'��MQ�g�4�1��e����i#�r��cks��{�����<ι�4�nw�(W����#;�[_�?�Q������9���"��fT��)��Y�K�>k�@��ɞx�{U�Nzr�GC��7��Ϳu`�s�+*������s ���k�;���d�[�e�F@�ų��ņ�Z!Pg�$b���
�a][�lSV;ƾ�R^&u�b��2ި-��L��d����|�m";I4[�]Ƅ4��[�ހ���PjAa��U7�PCSuӸb-�*��77'���e
��:y�?�oy5s�Rx�W�G!V�o�>!����9�v�� ���Mq�~��!��-ZubWB}⺙�������h^C�r��4������m��S�k��?2|+��1a�p���XK�iX�䎈O�.?�;�bQ��M���A�A����L}�es�lGGm�hm���������,��!��J�:�c��"c:�sv�c7k6l ���>��l�t��.�4��Q
����q3�-:��^!�p��d8Sa���B�Y-�ﳩ\k����̩I4�Vt�^�?��9��)��ބ��!������I#NBF����t�4z�z|ńr�|�	'@)��F��W����C@`&�)$���c­�6�${5���
����,��.q��� wu��a}^:P�	,��-F���r��D{#Eǖ���h[*�I'��sK���!��l��/�-no=�vc�48']��u[P�y�-Jw�n��*�y3 5e��Ŧ�7�|����|#[o0��SAa3������V�挮P�g���k�xIt��L������xɧ��t��ݩ��4�D>�T� ���`��v>b��0���Qc�q��$���8��u��/�(�0��@����ʫ�N��T��J�v�b� ��g�R9�q��,��� V~-SV+�b��l����h)�wWi�|��7'�	�Ř\�+���;�������������:��d�^�	 ���T�;_h����q���t�jg�O���u�O��)�$�w�%���jy|��Y#��T�����{���2�~��A�_j�3�(4��Û��+?�ݐ�CL� ޠ���ǣ=lPg��U1��{��}�'d3;(�u��i0��Y2��:�eM�x翗"��,���[gr��BeA����a�YT�W~�ܵx�rKj��3�@0{�?>|��*>F�ٮG.  �����]����[+T��O� S�\��I��rᶓ� ����h(���	Bʘz��-��d�;'/����N>����2pU;VHnz]׸L���۟"����h���@&��\^�{b2.0Co�廲w�Tw��t#>~�sa0�yІ̍�fjM�ԛ;���+�����ů{HZbfO�ل@�+�f��"[ck��^�;��J$'+�rS9�۽%�m&3yg^�G�����b��@-rV�s���d
�����h�Y_���^�O�WV0�!C�j�>`���;�B3��J�����_�Q�aƬ!ѽ���I�w�ҋ&b����As7[:�:�")Os��	��k�-�0w!Tre1�Q���H�/N0�d�{v��(��yw=���U}f�B�jg*�	ٹ,(�<aT�Q�S��\����th@Od5h�nF^�5r	m� �^�����d�,xv^��@GH��Y "\[��1ls�7���]'��D�{m�i.���Y=����B�=��췗%��堥֌���W��h��Ѩ�y^�EQ��߫`qQ�UWKn����r�2lŬ����.��"?�O��0jF?r-��e�K��y%SFA�b��`����8��?�|r��Ǯ�U��l�{ �R�����Z-�frܽ����32��F
>�r��>o�����n�i��[:#!�K��A�xriޱl�r`ӕ.�{rs��2d|&/�T�2T�*՟�Qm�%�k�^�=n��w
Yv��\#l�Ηۣl)�>}G���p"G�y�	 ��w�>���6x����J��L�ba���-�B8��;\�K�/]o�8�ja9S����u�����U�2d�&pS{|���?*�Zl�N��QA��&ظ���EƋG�#l��$�sS�y�W�-��0qF������,#��&�L���2\)dq9�{���!
j��/�*�E�UiU��ȷ������b6��D+S��޾����RƳ@��̪��ۖD�t<�a�O|������8]g��������}�G����t��4ј�'�@ݭm":("��8�������V���9@��_@( �u�gl"ю���/��<!�"���S��E
����{9H�n-�Md3S)}R�_�>�������O�Mxe��$�i\ QHto��)��8F�&J8Lu�^�1�s�3�c��np��q��nZ�h�K�N����cCY�"���<���3-կϰr0|fI�K�Z�ǲ�Ɉ-ڛR���`�?A���h�#�ҫ%�
Co�;�	jΙ��?b�}Z����X�� ��'���9ְ{=���ø
�@?wi��#��^�u���� ZQJ�S爰�JX�M��̗�ݸyKi�+��.�C ���Yp�9q��؋��@41b���#%$�쨍�$Y��g�M�8~���9w�[��G�?���}	Vv�f5��$YFő0�P��͘G�b���ʇ�1�Z���s��|�'�-�J.sZ/0i޹���Y[�.*�2����S���S���J�p�^v�l��r��4�CH�+nS�	�T�g�ƣ�Z����1����;����l-9��虛���3�x/S���\�*?�9�I�KYˠ���X�Y~m�悡ydϱp:M~:f�K�` M^�/�����\��[o�-�'
ղ�+3�$3��<;�IM"����٘�f�d��ubߘ^��n�����@�#���4��w�Ƃ@�׍�l�d!�˕0�	�v�M��z��Ţ�nV]�MU�&��ؒ�7I̽��[bl "7���	Ю7.4V�;�N�i�e��k�@���+�D�^3��՝�'Dzpbczn1Vk�"5�ں*xe��`a�8b���]l�o�j��I煁oW�(�E��am!A��s��Gw
�2�50"*�*�a� 3�.#�$�l3/3��, �A��WQ�s�y�˹�U��S����*��o�hl�~ ���JG"�cў��E���tXF�ն��h"bc���Ka�ت�î@���w*�e(t���XL�HV�n
^�=ݻ�y���`�Y �.�zA0q4t��j0"����F�� M���o�~�����������%@��A��xX�+�����b�f;+5I��w(�Q�
��՗��?"��Fhd9h���FTqU�G�6D43�����c�#K��-���:_, ���Vq<�W�H֘�9.o��/�rn�`�­9��Դ&����^���Z*t�G籥;��je%��|��(�X6 ����h�W��߃ޯPn���G5w�����֝v|alH��ل�f�'����&5�{���`ԎB�Z�n��|��Ź,(r�F@Ks|Sn�)W�2�#���{jRE��I���B��@򊙜��pQc͚��R����	�z�-�%8�z��LLl�5�Kr%(���P�U �S{�u}_�?#$�"+D7σ¥f�ǧMd�>C�y9�`i���0^�Kn��/�ʴU�pB$�Ly��q�����ʸ�]h��_��Lв�^2�@��x��w�R}c��?�x�JN�s�N�;�^%�d/��0]�i2�-��9/ �� ?���k�2L�v�cW/�jA�,��+�B�$��C�\A,#� J�-`$�n�7����'r|�iZ�f��H����B����3�9CD�`U�#CK��U!����%q�6/1�C ��fTˍG�zD�#��?+��Ɋ�8�N� ��`���!�k�P)�����v2�\�^Z]�%AqReю�� �`�I�~�3NKm/S#��w������!ۖ�{� Y����-T����/�	���[���1�G� ڡ�e�Z�jT�6RV��/��ì#kտ���Lde���{���������9���i�I�M�(�<y ��*�����X�[F�q0��ģ��zg3���Z�/�7�;�����*`K�j�O'߹9��E�9��G�Y��5k��O�O�Z1x�8��l°	��Z���{F��'�17��[T~�7#��膏9m��>.��K��TX�����E2Z�/���V�*�1�ޚ�<B\-e_r�����H��(OS�6�0��9n�Z�l����WK?��3Y#�m��=����0:��! w�Z�Ν�!�FJ[��*%���R�?�z
���oȰ�˝��K�~��>Or��B�t2�5���L�UIէ��= �H���ML�eB\��5)����� �0�2�\(.�J���0�5%��W	�xs���R�y3=��ϴ�͡�U{$��>n���񀾹`[�/
�5��E����'4�4�ҽ���8�P�n�Q���`;����/gj����!++%��m:��u�0.csx.�3�[�pR�߃1�LtO������X�y�@NX��Гo�dN#Q}v��V��eĆ48����9�$�miܖf�UEN(Ҁ��Qž�¦���MZ1�t��4�Me�Ws��b�K}r�㽁4O��Ke�ݣ�Y���z!�Y:Z�_D�5��z�� ��d%쾵I�Dٺ�`O��$y����oI��F�j"!�8v6�)pnZ>2-�I:���~���CF*�W�\M��&�%�y��B�U�.��:�8�V݅�[�*ć�F�f��5��WO����m��!4W������K�����&�z��'iQ{��\��Q�<��rO:��+��ɩ���>�-G��Z�%��N	Ԫ�
(��Yu0�˔U�bb#[��6��[�#t���y�����A���U��A_	��M����XY� fNT@z`W���c�%5��'s�77=2D�CU+>ssP.��)��:�W�$I����� �p7��(Yf9�rS+��V!?��Zp��κ��+�M_�bhg��Q��+3*��%范2�gA|+�����:��Q���6k����0����6ѥ��/�b�g�RD$�m�޷�yW5�'�%jc������&Êl��p|���������������;%8}8��O��,l�g^z뛱�:��7v��I����a�c߆�#>>��-�4��̳�Crj����.����7��sgM�8%�Qk����ͤ��i����|�����ҝ���DC����<M�j�A������t�6�Zg8ǣ^�xh�_F����ʖ�n��Q��C�sAh��Xǫ?�� �t�ˌ�J��w��F��"�!ʆbP�u�6x iIƓ��΃)�=�O���7�2f�)� ����!#�)T��1�
Z��c�a��֜$+j`�J	䓈#SP ��;�,ֻ� �KCNt�8�p�Q���%���9s\�>H�?Az3 ��8ut[�J������Ok0<��فf?Qd���* K��X��9[9���"麊`C ;�O�+w[1���Wqx�0��m:�k�����`U��¨�:q��-�{��v���eC@�/�]J衹6����y�u��Ӌ��z��m�g'J2��~��!���c:!�0$Z�Z�ػ���xQ�]�f�<�	��`�봕�����fz�'�Z7WD*Bs��UK�"Mj�ϦIl׺d mC�2�Q|w��fl�<"�+��Sy\K���rb�^/|h�e��'��M��"'`W��o	���ν�V��+�1"�O�w��I��jJ@�|��& ��� ���i k/�v���b���3佽�axZ���W��S/cǋ(a�~*S�1��ިR���)#�y>�7�f]�ўP�L6U2x+
@γi�/m[��ێ���T�{��j�� �X�y���?�]
2�d%���,�ہse0(���)¼F⻍�����y��@N-��S7<��4퓕�v�8hۀ����q�?��kP��td�{MhWh1���+��hU�@�]<1�@1S�J!���O�U���,�+V�#��F��'�]��|�JA�}4�XYȳ�#-�� �}��0yHE��!Y^�)�c�||�S?�`�^?� @�)�DF,�Y�\��6��a%:�=v�o�x��jA��4���.&�tBf�y�M��!�����K�z��u �d�}�X��?�~�qs��R�WA��0�fv%��R]k��Vn��螩P#2�#Iֆt|�۫������L��?a.�-T�_�o$.�&�
%h���Ѻ��h�/�� i�3�{-h�RK�d-a��Ո%�uB��]�f����u&s�`�W6(Zג�4ͦ�����/���3���f�s��΅s��gc��7MB���0�K���:d9?%Q9���x��x��z�Œ%e.Y��7P��.j$�W�L�I�6,�.��۱{��pr��n��Z���#sNۘ*(�ŗ���p!��}65�X�	��Lf����t�<�E6C��[v�LN�4I���z���jQw�q\�LE��N9A�0��T�O��cA�����(���X1n���ݸ/��䓃�I�JUuF��-����Q) K��1g�?�1'�wX��1��U�ڤa�o. ͜2�9k�1	Z��<��y���2�]v�
`�t��_l&n<�-�s��!���?z̖u>O�/��z~���k��@.4��YﮐK�G���~�8䷗U�D=�9����	ڪ����� ]ؕ-S�E�[�j%'���t�{��g;]����Z�-Ot	�z�'���`�]?�Y}�3y8EjE�f���T�^nSǅ7�u�H�:�b��̯wU-�J^�ȎGX�-@�2W��W��#�7-&~���1�/��������lx�"�D�)�w���J\ o�G�C�h��9�}��Tn]G�ʷ?�W������?��y�'r
H�aK4ԫ��A[�;JWK�m���+�Ut��a�|�-.�d�K5ړ���&	�$�ӣn��+Y隷�/�jҐ̒4�����(�uo}�azo�8:�U�_�S�e�'n<��	����:4���ζ���,J��4�ܭ�6���	8)g `�V*+�NW!q�=�f���jQ�v~�!gL�m��B��J���P��7\jr�C�3'�sF������Qr+x�ߪ& �# ivz^zq� ���q��v�'�Sn�{)n� ]����`mf�2G`s�N��(\�x.�&ǣZc�=AYU���.c(������aM����U���[�U���� ���M���4AP5����n*W(o��BE���L���ؙ�u�u�pjo�!<"h�RY�;*b�g��#uk�!���^N>P�]��2��_�컓V����߀�P��R�SI�h��	Y#���C1�����*�e������5)�˖��iY�o��q@3��M��:����������٣���_E�<�A���V��S�͑��"�ğ�2�a���cJnU�9'T��"�+�U�+��?K�l=`�Vzp��(	�+�C��9i���:��j��/���/:�Q7Z$!d��P�셮��պ��+ ���]M�^!����}a��w�Q1��|y�3\�:A���QI$hi����{v�\�\T���6u�Ac�hMiMU�i����q��6�S���p��u��˷Qx��z�m3|yU�p�{�~�k�Z��⋳�t�pH������_�ort�z�V
�����e=�}?��J����pϬ���~���~�h/�aSвؖ�ޚ#1΃�7��b�iѢ͸P}���X{�n|Nq~����ؓ��9@��Pi���%^J�V̷(�c��l+�ķ�M#��6���~�y� ��j��%����Q_³֑E~�,�6'1�!���|�'L��k1r�
Z+�9���Z��D�<�=�$�Y,upϐb�R.�""��Y[/H(�+����N��4o���r_vA /��~Z��e�N2�p����g�a�4�_�1M�u,��a��!��q��-6[�D+��Q��S�,�bB�6>+$� 6@Mߜ1���ܓ�p~V1c�CT�p]��T#���G��Q�.��.��L~)
Sx@$VG��.GV�~���+1s�*��.�i%�ۏ�5� u�GGh�����NQ�/�^�AnA)}��؈���O����d���y�\�uʞl��,
�RQ��U���Sf3�O�b��{U����D;r��a��w죟/-�S��1�?��Sy&w�ۭ��B��U)�P�A��DJ�a
_G���N����Y��6��#uCD��QP������]:��ǎ�oh�%�b�L��
'`#�6�ϸSH��҆H��_�X��+���B��\�m�\O���I{Q)�l�D����R6dޡ�h=NXܤy�~���v����js��79|�\g�Ar�������p�N7$s�F��^�#�O����>� ��f��C	G���=�k	OƠ�2�)f������|�4��l!ݩ>p�5u��������FK�;E@��S������t4�=��ӼG��Z4�B�X�u�jk������f��F|h���͜~ �c4��8�B��P��<nF�hjX���f�z��8�5�pDiUN�0s)D�I`��_O��3��;�/��;m|��-��G4�x���ʯ�P��G �r�:0yRQ��[͊����P䋭���Ę��p�2��V�(�<���fr�RZ�p�M���c�'���M��� ���k]0��0x�%���K����mz�ȕΥ����.�L�R���"Y�"p/����â�����-��K'��+o�lx�\;��\}g>��)=����Fj��T����� 2m[�l&�3�C��W�Q8m�����1����:y������%9؍���b>�4�y�b���W�[ė��W���3/��6� ����Z��^�vas�������OҶ�~6E�G{��*P_	��j�M��8�Nތ�6_���nP��%?��x���%)�V�攧�%f��]�.��.����ڋ�������Px;lL���w~��b�V)�Ո� v��dף�0+�-O��5��9wx܋�yj,�w0A��S��fp#�v/Ks~aSM �w��P#4�˞G�X���6t*6��q�RR�obS�hu4_\����X
X�#�6��;ޞu��arػHĭ�}P���dx۞U�Y΂�����l��!����ܘ�d�p��X��L}Z�Z��H^�T/)k��K� �pO'9����Q2_������q_�{|y|�Q��G��(�������)��H]�����Q?��>y��~��]H���F6*	4��֖��dz���#��B��PZ?�8�Ipf�����R�ǲr�s�ߋ���Q%��K	��G(�����BK�9��rZ �	=�5���u��0��Ң˟�L�J� վPD��h�>���ߴ�!�/4�� &�U{�
��P~Z�r�*��{�DM�����jMRh�h�2�:���Ƚү%]����]��P��Zo�(A�D�a����IQ5K��b�OY<0=�+�8�3�y�}�Mr�^Ֆy���8�MX-��?V���fdD�Cmq�CD-������I������+�x�i�_X������$��D��׋�)�UuIA݁��2$�� �h滯��_wc8�������F��b�l��^B1u��Ʉ1S���V:�T�s�#oXQ���qn$�������$Ͼ*�T��g��}��R�ҙd�<D�ӳ�ڵ��K@Oy�@T��HP�f��bwm �,��F��&�K�����|�"x���� 5_3�ё����]�hZԀ�R��w�)|TL�F�v�i�X�k8�02����;^��,�@�����z��H�nfR�����e-i2̡zH��∁�w��/,�ēk���^]��RR���� �	̞̱N���VἘdYg�%yߕ�َW��X��o$B��Np׿h�?Yz��y�a�UW�iQ��RGA��X�K��`㘸\��{p�qef� �.���6�,�����-�+:�{�N�P;=`��=]���r}�����hf��Ey��l�����C��I����w���
>WFVaL6�9~u�Kk��E6�族qͬx���A�[�<Gh%ښG�,^��/}X��lО,2��qμ�z2n �Ao8j9�\������t���0���A�?-�ofe��|Z�H����9�y�(�EE�?���@Ɗߛp��vP��i� �	�Ǉ�Z�k�?Vm������v��>��t�a���k��d�>[�E�"bA0$�r��"�r��[��)�W��t���� ƭ�0b��D���T�-0���l5��X8���J��it0k:�t7�wu�2���=����W�v��8�t17��bFI�C]�^`�#�I�S�+��6;���$)bj-���N����^��[7ԲC[uu����%�<;�<��l�1�.D1_�L<i3�����Y5Mog��ٴQG�0���è�(_���J�ZC�u�PE���Ӥ��?�����e�]�u�Zn=��Q��P�8\˟)��.�s�Q�4��o�Һ��Z���c�+V,�7��L����lV��.L��s�.ѯ���	��JGe\�/]tP�����)-�= e������ܿ2��d֓�m���k��×�J_ꊰ���K%R�k�M�gk�m[����a�P"����Pkeˁy�c�oe��.��G����	�r|�7}) GZs:z�[�}�������U�Wl�-��0���u����L�����~��wI�'<Ѫ*R�����k�-t�jѬ2�����Z텑]_���(��)�t�<9�q��;��i���6���C�W�ڔh�$Z�󶶵�^ߖ����g��=ΙI������[o��2j�	�t��(
�Nw74Yߞ��O�Զ�!e��0y����9@���)q�����V�~!n��3,��rq)�����O��9����%C��£a��F��������m�&I�D�uv	+f6�dĖ����e��GЂ���2�r���y.1��y]�T����*�?��Qs���E>���H,�T$����|s݃"�Y�E�-�	u�fU"_�2�[�p�lZ��y̌�K�nF��y����}R����k
�qԉK��}�@��W�N���aS�ӑ����S��8~��*~j���Ž؜j�U�9ޅ1��Mkث�dQ����<��`p��p�H�WE-U
,�FГ\��r���L"��k��|5�a�e'2�*J[��;�%c/�U�_�D�z���?�=wL���t.XH���KHa��`F�(�].˾�S1N}���~�Q�l��|��C'�����`G�{��-o�Fh5��H;\�ö̽���*�� ��QG��3�02g���uD"�P���X?�{��Hh�e��ݢ���:A�����Tp�bz]:����@���^�YQ ��L.�t����9�^ȟ³�i�����K	���UU����BC���iv���5�SW� ����(�o�ĝ�ic`�9n{1"��·�����]%�&m�?Y6����,���|]U �Ma퀜����/��L����[�3L�J*���Y�ں�]���]�z"֑۽�d��5��ċX3�q��,Ѷ���8��:'<�0;�����{o���mMj?���V.sKl�F�5�$�Y�Za�%�<KxS����)RFsӍ��c����I.��G2��[��D���,@��C%���F�3�~$} K S�~>����6��=ޘ6�?kS8;,G������zv� �q��?G=�P�4-D��#>STNÜ�u�Ta���E��"&�#|gD���H"M�(Kme?Ћ4X�����aWw�-*�l+������t��<Ϗ�cۥ	���7u��Q�F��!,4�fҏ|L@�;�Gى�ˢ�RjE#��朁.0d)'�r�)Z��� z�0D؆��)o�_�h2��+�Ť�f�X��1�o�ʀC�B��WAZ�'����2S�O�J��G=Ϸk�%p�!���2Ŕ���*g�7�](mu�A�g�Eg/c	�G�0�[<��	�G+`����|���/�,IМ�z��m��T��]���[�$3G�V��XP�b1=�2��ѲZ����ҥ��%�;����]�.������׆���ou���L
<���L&�$
�>V�w橃?m0i���-|y�p��=�JA�E�wH��c���*U��7l9�z�|�b�W}�s�&��9��Z��(&�T��"�b%{�4�R._��E�R;�W����~K�".�c�e<�-=����i�ݱB�B�8�^�D	��.t�g�E6R��7���������TL&���o��O��/�F�7��������6�C,L8���I��ծ�
���4Uc�!��6k�t��V�P�ŝd�YN5C89�z
C ����QT�Ԥ�4ny�Lp�� f1BŖ�ͫ�̖*׉p�$<�+Z�djf����/�Q7'��P���6f���C�pP�u�"��=�Y����i���ل_��^�Zlk�X�h:�q'�C��ٚà�������=�u�ǊR��N��l1g���tf&J�K`ʹ��������﨎 �]#�D���V�7	z�p�-��������=R�T�}
S�EU�6qT�d��m6Q�w����9�M�Q�wD�zp�g�o*��c��oE�Cy����o>������s�O��>eU`?Ų
�t�{V���� ��'�����9k�I�f�TA�U�����n�Z�_J���$!�ob��n�dԾSa�y����%`b��7��Zx:�� i����^��h�e�eW���zC<E]���Yۢ#uZ=j7�U����0�SN��Ѭ�f���$s�#W���7ZMAF�x����p��$��_���f�a�N���/�;L(j�~<2	9zŉB�w�
@}����W���yA(��@�C��!ICs8��t���g���z�Ĉ��p���fx�&�?�QJ,Y�!������5�f��3����>�J�
j���9��}��n.\���z���pG���c��ݕ<I�)E7��@�C�v�Tu��������2^���X%��Zy��E�+�����=4f��x��0HN�Zt_�J�hy.��i��jJ{�[����luBN�+sr��i����C�Ǚ��r ��� ��@(�&�1���`~�\�,pVE4�˷V�`�V�|*���Oܻ����?�'���k�r�q1ȁ���B�k��U|��c�?`ʕ��&��\~���3����a�|Y@Yd�WNәp�c��lwa��'��l�%S�w5�$��s�#048����YD��;]K�A���8s�"��?Db����=Ē�=�!�ϙN����J��6�#����/��w��!y�x*�R��#�Q�R���o^e���]�|�
9r�Yۜ�� �7�@��NG�cZ��ʜ�k>h{r�;&�Gר���n�Cx�%�>	�@�Pm��%KWA,����zOZN?������X̻�Ast�/Ӯ0��u�	�$녳�e��w�T��o!���xUh�xE�$sʪ00��0=c��f��SZE5�3b��֌Q���@!�-I�n&��I5��f���2�m�/i���|=�A��ԗ�����E(��(#i�cYY��:����Cf��ge�O�y&�������hJ�*���+�l��d��.0��F8.�f�N�S/�_��>W9NȰ�{]�B5�]�Z����`�*y���+n��|�
Zc�=�w󰍹�&� �����4�Z�f撠�a��� �n��ʸ��P{y�7V�p���c�ݔJ�������6��n�F����f�^ߩ�@2��o������i#a;t���j�nvB���ցk0�F�S[��վ�)-/��0?��d\6S�Xq[F2n�b�0ax~���Ě�DZ��Dz����J��iZ[���&ϯ��MbV����,��ĺLغ��0R�g�آ
	�̣ɑ S�yd`��2c?z�KH Ȅ�U���3h������y�=)'�n�DF0�!���_�3��4��9d��(�J:��C���EL���q<��(9S3����Z��՚ �h�F��x���lb�z�T�`���W�)�%cjO�
qq�W��#w�J�Q�_���?�5�i�t�i�%����,��/���y�=���$.�����������h��m
d�5��c���^zX��T��D�Fj_�ӯ�!�����ٍپ7���
:d���>���V�G�R�g�mR"��b��u?o��eЪ\Ǆz$j�_�
��|���^�Rʜ?m���#�ҭXx�#OjO�n8ۊ�b_� ��hFH:�4�T�j}iyh��*&���֊�t��P"�/V:�6�9�QD(�Úm�@��t�&������6���I��;�\�{l��S���.r�F
�[�i��p>���ȧ����F�lL�C�8i�lW�3�8PP��&�jq�s�
}�R��?����$��`�Y��R��\m0D
���U?g>5Bu�=BJ/��E[!\Ġghx��-2���]�����ҍ��N�<Mbk)uz��l����]���D#Z�bz�h֐�yS@�MX#�T�b�ⱷ ����ə�@5D���s�p��C3�������:�gciW���]����BJ�*ѼB۸q�C�O!�w�;�L��R�]@.a:t 1>�n�WL����v����~��7����S;mp�
K���\��hc�O���>�<�jYh�`�
3߫�cK:*���xsz�IA<��ᇵ򑰅=
��[�w�ovF�恨�N��v۪-+�����S@��sj�~ɼ��J�d֥�p��a�����b�.!�L��;6��U(q,�t�vǄ5\�
 E^�9D�S�~f�OqǊ��|٥�Co�6.`�e�h���?����%�@�<� fՍ�@K�Gk��p��
$�vU�+����~
��������z���)��Jd�N��II?�ط7?Q\�o�OMΜ�Ý�͓yz1k��	�:x���:V@�MYD[�]/J��/�Kh�S��_��@x����s��C��>�i��}�,v,.�Sn_����`s]=<6��>�Ɣ�J�3�!n�[��\
a���O�E��䨋�H{�L����~��ˇG����x�O�PA�(),/���b)�\�-�
�0�j!]�.&".����"��A*�i�D̪�f@l��/3��>���s��댎_�?���Z�иm;�h�9V[��a�J�}C+��H�SK��c2RM�0� ��װZ}��p�t#����ϱ�`o�zA�n�3�$��4��&%��O^�8�pl��2���P�oD'��3ؚ��M$��-H=�`�)3��Ľ����`��U�!G�g�>�yr���~���2���M�k��;a�9��d��v���q;�#G��yc�h��v��$���D�.��PNPIwQ�Y�+�f"�\�&3�5%9�ԎuH�'� ;�q�F�^�7"�O�B���Z)9�5� ���\��S?-.�M�a����?j��̎duM<�bYp��.����r��]e̥�RZ:v�?�?��kZ�_�)
ueA���0?0E�u�^W`G)��%�yX�9L!3*���u�0�N6$&�$N]���nǇ~g'�~L���z+��xC���#7�G����:�/*ܗ����o��])�i^O��ؘy�Y���a�B��S"�)�L�.���HC�;�ka�mm����Ѧް��U��8�|��y��@f"b�����Z\˜�R�%y���H�_����9Y��P��O��C�X������9ϒ*�?��#&�ٗ���x-�|�i5ۀ�70m�v��d���fD��T���t�М�㳄��K�����Rs&������S�}���i�>:��ui�گ�ȳ�@���;�''y�6E�����Qt��)4�b*M:�v�2nӄ3����A3���Ȳe�vn�L�����ɹ~��>(�ϡ��9R{A���ֻ@N�'�8�e�3�ݐ��,D��ӄ؇"�I�0fڧe�L]�ffH
�X��DM/��#ŭ*�6�fͨü9�EU�Y<�o5�Ԃ<~<�H�f:�a��岾��֜�o�|� i�t�0�p���-$�M��oʉ��P�K��Zo2&Ɍ�QN�k�c�M�ԝ�'/��^l7$JӚ��Q��Z#��Ie������˭:��� �n.)f��d�>�LԈ���U���T���湥�n�@�;�����B����?�/B�$(�u���[��O�ˁ$��a������ U���&	��b�P��xuv���q@,[���i|=G'��Sp8��Â�E3 #�����%�KrP�����#���ܗ�j��%���U�
$�V���IIh��⌁? =d�hz;��X+S�~b�PX�$�J`Ĝ���m�V}/4(KqH���^;J���7&R{18���l���iD���
|5馸�_J��*#x�/))ܦ�f�	(R���yhzL��4�4]3}2�LJU3�w��[j�i�h��u&�V��`Y�d;k��� _�\��]O�#��$G�}O%{�Pb���d	ۜz���Ţ��ٗ�S���YQ�~���[\j;�0dk¿'�kK\f^�zㄵ�6�H;�׶�Wz^H,�J�'�c���~҄/��P�HG��Ϸ��-�ڕ����+9��vS�~S{}�	��ddR$=��J:�H�n Y�Ճv�ר6�y$�XĄ��_�ܤ���C�9��O�\��W:W8��XG����?�����������wߜ���T�ec���ڭ�g`�(sP��X<�&��=�-[2u���V뿩��-�gWx���j�����i�c���0f�*��h�&�]�&(����$��7=گ���{47��������aP��Of�H%�h�A���ѝ���Pc6	��TM�0L��Y��c�������h2k�h/Ӗ�X��c��IS"�ς�k�g����QqL|˿�fWJu�!��"��(C��1�S�"Uw�8FOPD�Xr�^Ga��R,�}���v��� 00�{P��k���0+L���56���
݀�^��0�K[8��!�v��uYs<j�&�R���^�6�e�Yz�Uh�I�Ca�2N�S�" �C+@w^.s�F�נq.��[�����wo:���zc����̰#o�@KPOw����~�ڋX�xH A`��j����L�����`����	�M܃���uԭGBAk�>$�[>[r����^h-'V�k���U�(	�,k+�D�e�\�I�noo�?Fj�c����ë�@��_NY,m䈓a?ʰ���	�lsD��f�p����U�R���L�����qZ٪���b�jL��{͖��ۭ�`���5��h�{E6L,x6!�2�[Wa�F(�1�����EE���G���OU��1�I#�Fޱ@�|�B˒�]�(�>r���G!~E}�0��K�u��'U��6�M��
�-�O���T~�h��H�{1u�����ZzI��,VD��q���Z-]�ޗ.��v�t�(v�z��wΰS?)�[���x��;"�O�����������q�~]�d��+P�.�"�����./�g�Y(<0�LOb��.9s;��f�g�^p�ِ*�kU�界��n������a��(Wq_���A79*y��&�n�����H�뻈%J��5�|`�*�zݥ�[�``����G��%;4�ʜ2v6�J�Ȧ�
� 4�<���ǹ? �g����9|u��=�|�N|>Z�FS��u":]�0F�:��Mㅱ�� ��.\�n�-�,�$l�����d��IaQ�ɋ�)�^u�|<�UY��H@QCUphp�xj��=霴'��zy)��l�q(�L#k7i�+W[	m�H.��I��jG�|�%�Wum)���&��@=e"�f�fk�$��W��B�z��ao����f�ӘB ��?��N)���ҘVa#���4�a�F?�r��5�y�������0y�R��{`�G������
U��q�g?��TC[Ǝ=��Q�qn&�j�E.��d��L�VÐ��.���� Q� � +aq����C�y�f1��R: R�h�_S�x�x]��S���̍̓%B^�o�'�^	!�'���qK�>������v�ff�3��g�2aL�49��4_Is��i��xv�>�_�N��sr)�D�S�]�+_=l8�)�:N���i.��|��2���cT/s\-z58M�[��p*ؚoI��~�a^�z:x�ܩ��LN�����g�� ɡA��QW�ø�R�߯�_ӄW�Q�Pb�������c�3f܄���L5��b�:W;	B�����/SV�NQ[�繘�>ގ�&{��������kQrJ�U!xy	~�bKi�_�,�:���F}��נ���k�q����*����T[k4�L�bSw��3�ݡ��)e�@�7�ɶJ�DV44����x4��G��g�1n�ºӫr�z!0��UИ�clW|�����yIӝC�eQqU�t���baed��P�f�dj�2��g��M�x�"d;Ʒ�,��1�W��{�l52�+��4r��'ܜ��L25� ����R�����Z\;�>TdY���9�jh~�M��b��R�KG�W���[� ͨM7/7��t1��b:�~����r�T�h�}P��n�] �Z��p��.8+Ӂ0�O�E�<f!F�Y6 ٢]��(fn�a�F�x�ԕm�^�ׯ,�y����-1�[$��3@X��Ќ"�j��C:i�#|h�Εc�t�l-S3w��'�5t��I��D�Ǳ����<{��E�	�[3��A�������H�ņI�޹]ؐp�J5O�u�5R��k����cJ�%�CW�ăc��	�P�3�h��"^hl��e�voP�����-�tAu��lk���M��I@�9d��iȠ���^C��X�6�H`�F��v�`��#,8��n!�����2�}�> ��<!9*��/*����<I��T� ���5�yR�]N4�N�
��[r�>b�l� a�z3?k�I�.o��F8��L�6��\�bk�1t���'�{y���+����1y�@���OJ�/�,N�!�QD���4К���C���+�j<���H	��{�Î��8O�L��-.��� �K��]�m�>��r2�U�h ߅G-m�bX����eZn	�I��,��WF&��# ֟��#v1��T# z�>Us�ZL"��c��/ֻ+)�Mp���i�Pp��
B�f�t}]i(C�Q���l�����U��ջ^�D�i5���^7��Y��!yXGB=������~'��#�6�?B3�VQ�	�
bݴs��Q�
�kN�,#tͦ�bEj��*�Ţ3f5�Z�3�FK����o��*eM�d�[|B-����~b�?h�F�8pA�];p�y2��ρs�x��823�O�<�*���,$+�\t�%��{���N�٣����-�l<9�w|cki��
��KF��	��k.�zW���k-�{�ao��*�]�,�W7��2Pwۊ���:3y�]���r<$��k��"K�YمWrm���^X�9TĮ��0�n�G�����E�� 7D]f#�7��cq��'�-�Y�D�56)��;߭1�d��4��s
ͅ�(���Z6���L����zD�H�����$�9WR{;�!�^��c��`��|\��ce���ts\
�D`�xur�,h��`y�T��ƨzO���o�mLZ���޷��N��%��NkX���!���r3G���5�F��{��56>&�	�E�k�M��ªE��y�f|b�h���`bC��W(Avі{�{��]�#��8��d�e�P�{��/�E��°Ȝ��}�i���$�̘�a���-1���)�g������;gI��"2�}@��P�\�t�T~�����UgFב+\EϠ������Rm�{R���ԭj���.F%\�O.�bd�iDqI�_��G:�Q���ʬmwsʱ ;�cI�B�yF��(�Zzo��p���h(Q�	�*B1w�|���A� .M/m����}�:>9a8�WU̸�6G �u% �xk�+�{����t��O��|;Q�<��C	}����&���L�ƿ�9����j�T�:w��&{�j���f",��,vΗ�҈�3JL��Q��$m]l��M�V�8kM�ڔ��׶�b�m���"6�*N> �P8Ձ(X��r+>S���e<�1��^�ԅDn�5�9�>����������A�Ǡ��wn��j�t�s^�m!����޵ަe���})"`�NA�T���]O@x���j
�`7bR�iK��#�TӱVŋ��w��Y3�C�=��+*A���*j�����x�B\��MX��i`�9�A���~��V� z�9�����)v��n�".�_1f:����5���h�-J�|xF瘡=E
���'� ��[Z��[|E��T<��F�jq�W�<�8Ou��@��
yJ.���c���OU+����-a�]4xC}���^��B���SP	ˍ�skV.�M�#\z�  A׋��=>3�[�М4�#UcR�)y-���m
��a� �
�¬-886��� �N<����MQ<�jv�iY(�w�8p�����)�YR9E=;�vn31���:C~�U�L��4�v\����#]���:�o%�T��A
^0��$r>��t�LΘzȱٵD^�v-U��V�W]���:A(3�bY��}��baI����Uc]�3���y�@k#ˌ�-o�[QƮ7�<�L�42m�z|c�
�H<�����؅�(����b��˜�M!��Maj���w����`�/8s�H�a슋q��B���2����{�({�G
Qꫢ��>�̑�n��:z�p�I@	ξ��a"�)�����%�w�PV��E��^�#j�yObz^�m��U�<�|��HO �J,��k�/���*����H�d�����ȷ��D8�X>n�H�qg�S��S*8P؊!R7�+��4��f��!�
�Z<K��H��ղG��(%����.S
�6)w�>D�� 8Q��H�C�lBGu9�b/�Q���A��͑TQ�3�P/J�;P�[�V�C+ldI拿J��%#�?����Nb����sLe���2�1�}�C�㢹��"��d����hfZ�~;}��V���|%j}���� 윰3�}; ��!�0/�WFQQ� �*$5somK���x��o$�<wb nsK�0�0��\21�c)�a#�G2㟛8K�0��@8zj��N�G�:N�ܕ�T���?�/5�$}� ����Cqx*;#`�gfl��_n:i���۝�R[���I*�~�ŗ���[����0x�f����p�~��W��V0����;whV-�~hǧ�
l�HD����!L�{��fx҉����#�]��v�޹�q���/���K}�b�U|��-v� ՘�ebz�_s=g%�h�o�\kW��`��#���u�t188t��;2���$}�jQJ��2,3�rY�\0��h=�$`�U�*؈�~v������jJ=��`a4�IdL�V�͸G=W�f�g}h�6��ye[�,oA�� ���Ő�5g�E:�)�gc��܉�t��A�PMt���>���9����wA�>�c���Ҥm�n;��!`eK�;z�s���7,(�^�I U�����p� ��RZ��lH���E+�?�xfL$�s3�Utq��*�FnY���R6[eX����4j�8	47��$4>�tSB�����jǯR\��c�i�\��⽶�0[*;��E�����\��0��mZ���ΓT��KXť�H~���uê��x���ԃ����������w�du
s=8b*�$=,Rb���gT1F�Q�x�+A�����c%�+��B6pK�̔�a����$�_2���)\,F!юY"��NÜs��ݞ�]� ��8��x��k�t%���3�؊�H��q���rV]��z�j`u��;�B�l�����ﳞ"���o�Xx���/�+�\x;�q�����̅X�+Ff^��]+N^����ƌ�ކ��_�:��L��TV?�J
�������t�C���Q�=o~��j�Эc^�ʼ�9b��Ɂ�[� ���+*���2.`W���)��[\�i�4�Q\���?(Ȏ�߽����a�f�Q�"V�b��J���lE]a��᪖�2�U~����@7���Ql�7�i<��wi�R���]�pI���*hT��T�盼�W��%@��{wn~��5B;l���5P��7�tGڀ����gњ��b��c����;}�������8;�8�h�	o}ͼ02��"�$�tC<�Al�l������D� >l�u'�d@�7R��8�(����C����iMq����	�O�[3�@%�L�@0'"��:m �Ԡ[�VUH\��(��1�1����[�8�|嘸ZQ��T�&K���q��0j�״@�V��!�
D�rͦ��l�~���Sʹ�|����1�Wh�0*��v
D�>~^�2��qEq{����/����|9p?����WD��7893��RR�����@�>�f��
_1�vV�p��NS�w��?z�ݐ[��5�=O����|����
y+���O�qf�S����rߔ�<��*
Ӷ�V��E�e�uH��# ��8���G���F��֍��^E�+��
����B�K�r�i�%ѥ�te	���n�nk݂,~_W2*�"�[�(�`�Xчہ~���;�x.�H{�T��5�������e����6X�3�{��c6�u�/�S|�/�G�G�~`Eux�3�CsUzxؙ��9Ӣ��Q���@��s0L�^�|I����ݦv�*���L�Y�i1W�<���5�X5'��}t
9@%��ӌ�ٷ3uLr!��&<_�6����
4��V���qI�z���O��t4�K+(�X�ۀ��|�B�d0ܸ�w����@�?�;�͡�@�������3c~>7�F�"J�3�R'
��Nfo|�U]��nJ�~L)���kY�m�S��b�m�0�ڛQ\��d�R!@�5��� ��`�����&�f��Y�y�d��M�Ae�5��c��Pم ?H*��w���q��&Sm���f�b�wu�n��D��(��1�&*��u���,�[� �W�L�+h�.0��\v�d������
�GR�n���%t�Ҹ���<�Pc���怠�!I%�gKG��}�ʂ�:X���ΨeÅ��q)uG�:��hl���o3�����آ%s�|�;�i[� Ao=�h7��
�f��ß�4];�Q�<دk�����J�(A�P�&�#�1ӧL�����M�y#��{r���[w9��	J�ca�"��YFE΂Y V#�������L@�u�펾m��؄�
C��G'��;C�Z�UEZ�­��m�7�5XY���`����y�o�-�I?������Ef'/��29����Gt�'brp˞��e�p��.N{�R���]8>�_�=��E�2 I�c�ȉ�B�XNf�(;0s�=���gk�������F�r<��#�Ϛ���q���e���}�bݓiQ��&������;�/�M���=��*,�"��<J�e�q���:獪.����P��.�y6�0~��3���������Ll���U*�g�m�m��݈�ICo����[��BX�o0 �>���A�A�'�����=�dw �S+��㊐��QV��ҦIݼ�����AU�@�_1�ՆJe�<3��w�Tжb�FKd�E�׭A���D��~Tc���ۦEq�,	ߗ�CC~��r���O��뇟�y�T�j`Ů��cZ�(��u�Q�G��0������mWA��!3}Ծ�Z^`?d�]�{v��]�s���Qy��WAS4�Z۟�5CDV�����_ݍBk����q]�L�;��O�R#�#~�m+,�i�Է	DO�����%�*��)��nT�D�9��qN��~Mn���!��y:�:IR��c=ܘD�E\mIj!{���
�{P�`D��{���~�>��v���2c$I�!�>�"�ó�Ma�݆y��*�sXz�AEB!oVx"g �Ua���E�C<t��"�K�M������63��#:bSB]ݛ��w߼W��W&�R����rX~�������ǫ�+����*����Ԕ1;�}P쎡	�E�j^��g�.��<<(�3�����`�~b��9�f�E�c5dߛ��hoK�0W�.�[��<��E��bG�ZvM����
���HW�OBdu���݋�a�?���ڛ�K�M\9RG����(�H8_-�5�>r:b3O�tq����12�[�o��q̙�sU�L���$죴��#�t�+z�XP�T�i̮A^���y�f������9<-%$��!��<�t�
q��=�&��[��-�E6	����=��V.�[�@K�*�^e��s����.�J�X��<���ʘ(�01�ߢ�^��5�i����<RPY��y]�'!����df>�Qv���`�%��W������QÆ�(���9���<9����t��C�yL�a���b5��k�@����͌v��� Ka��ʖoǸMP����V�0�	h��4�M�*e�6e>�=�PV\pm�AyN!������gkvA�h�?��~�ſ.B�a ������q�ڶ
Į�͞�Wʨʡu���۵ѠǶn�f@J�{�Jh ��"����< �|���kG�͏X�oƋ}Kz�V��7��}�q �%	_�� P��t<����+�QP��rVH�|AH>��]Pܤ�-���i��1���:���ǭy�@}z������;���M3�:����,����?��.���A�w�����- �$o��Ն��5��f���P�G ��?z��deZm$txc�n��}��{�n�c|�Q�867pƘ@�?_|ɉ�U�.��@��p:����ҭ(��0Ԥdg�������YI�2���w-cFF�na:�gx�P����Gg�����b��w��}��V�Խ����;(rc8�U����Ŵ�X4fg	��tZƦ�^����a߻w*�Hߓ3w��ԍ�����z_Vr#����&5i�X<�Ȣjzf=`����:��3�\�{M㬥�����%\h����+�<�`��}����=�R_��(�Q@��H*�ߒ�b_wGʩ�R��)�
BV�f.��w
�VXBT<��5����[�Ň�U�ж/ z�|d�<X[;}�a���1L�is��`��0���&���!1&Ô�j��/ʺ:BS�� B��]b��
�u5��Ğd���3׬�������*9k	��|w��K��ƒ�,�+�1�rҤ:���ϭ���נ��ё�0�_���ݚ�N���b��'g�g��筦@ix���g�¨��h���n��m�a�ʱ�c|y�RA&P�r1�q�dM�є\o�fK]a�3?�8����5�+0e�����`����H�.g�"�wY��A���Q-�@-����g5���V9��Z���(�)%��iVkʛ�F{���A��S��98�cJ]���u,4~˪Ti�߆ӎ^�I�[tz��z �<�Z�`ݠa�x��LRY���2�xfFq����)8���0��R>��n���}��/������G�g�9`�Ψ��Rـ��XС9g����D]ZL���M�{G��4�������p����C����a�ʿʚ?����t�}�-a�Л�)�$�4��G�%��,����ǵ��Ny���>(k����ob$JHҍ<0ZZ��<	F"#J���m������˞҇9>�8/ρ$'��/�NA�'������m1���P�7����wҋ�O��a��G�WY��5d�j@,�����<�<W	<B�������W(�5t�(3�*W|���~�_���¼���RE�˺%��5�r�/�'z�|�w���!�J���2��j��A�(�5�i���<��:E���lE��bw��U=6y�t�^��m�����ߨ���~��j�q�E��1��{�ְy�Ǝ�[Xt	P|����m84�R?������wz�Yӯ��l*C�<ki/�1f����,�C��,$��Cֺ,g�kc.�Ȭz\�^Z}<� �S*�r�q�7"}���V,=[b�]c�`�3��vE������������l;Ao�#z���������[��g&�Vy�r�%�*�2�=�u���uܽS'Y	m �R|�!pａ�ׄ�]�oEeMo*�,6��>�WJZ�v��d������[x�\�(��?槄y��9�}��3.r ��VZ��U�����%����g?�e��A��%�2�o�z��J�} �?x�J=�ɀ9��vq���W���`Ȓ�~#�W00c[	I�#(G����)_Y4g�p'��^&΢�Ja};�AF�Y�ӑ�b�B���yfݖy�Z
�)��o�
t�;�x�wН&�6.��gV"<��;�ȹ�^�炌8��g�M���x���I<R�{�%ێ�$���,N���6;�e6i=���;��Am�F*��6���׺ei]��3P��s<{VQƮ9��y8"�`��	�m<�zlt�F�>�������Vܯ*m<g������y����|�&�'�&��k��Ly�4��h�I��0��'o%a�sv�T���@���24�=�I~�/��d
�s!S��ͩv[�� ���rq|Q�+I�
�,��5��K|c�*�Y�X�zp��xc��� �>��0�4���w��d\��m���c�����7�e
V���h�w�zJ�QX��׆����W�9�a�}�u��J� ��� �!�H�7��%F�+iP�m����k�U�~���/+_���@y��M��3J��z���H�erg¡���h̢ �8��}���Y"��u�*Yg����	0��k�ml~�)k2G}`��u���a�a�?�p��4�� �%�����%���z$E���0t��D�s�9���t�D��[�9&�3���hQ��^��Z��f�W��P6�%�v#�q�s���
���:q�2yr?�v(b{����no��STcy~�7{&U����Ap~��<��Mb~�'�+;����z��spP��\�o��,�],@�[�����_i�N�� �2�����>����+��S���Tc��G��O�ؔ����G��x����{#A4�Gs'֟���%��ÿgj�H-�����k ��%.�c�p���:���7����C����^�a[�P��D���reS����X��x��$E]8�<<},���u8֟f�1��Z���y�S��n��_��l0�ŉm��<��� N�S�~�p}�r��DÁ�f��}�՗�&#��=�n@���.�����r�aĢ!�����8�N�c���(��W��^>�o��g����sH� �ᓌnfɓ����h��h�������
o}0�۳�����FX�!��&AI h���aO���rr
C�����R}���l��;<�df�3�ŀ8� {�k� I$[�#Mط<�Q4H��53�bރG����o��K��Ӷ�Ҧ��$w�O��ۻf���3����Y+s>��+��`C�Wڹ�~�Y���ֳk�$��$x�EZn�Wv�ҝ��*��bH9Ԣ�u��xz�[�g��.h�zm��!�Pr2F{�!�Bz�t�m�o-�[�[$qkMb:)� �!#Y	����w
\�-�I��\5g�L�W$��vx�-�������g���D� �����s�,ٿPo�{ϖ�٩�{�?\��v,1R̀G؊��g��%�GX���@[1��J{G�y��),���^*�
��@��b�Wf�c��-z���*ػ�]�~������oKUHXH�6\]OcAe�#��ʗ��=6�#dY2����s�g�d�L��?��-!u-k� u������ �'��7�[2����_(��7��lo�R���VU����o�8���kza�-�N@9��B	�CcL���<Uܞg����Bd��@�`����n�U��@
q��>�8#��BQY	�_��t"$��+����K6�he�� E����z����\�<�Y��	�Bz�QYP�?���\_�����鿿>�_̇ϕC��@v��6��{]���h�m�럟=����@��d� �����PF}z-eT�߮_��{Q�u�9��'�jʯ����$�%B���F:�-G� �%��ּ�$7W���e8~���͹G���,��&	�N��y��R2�!`�,��Q����&n�h˿�\�:?x��l����]���rG� L=c(O�Bf|N�b�CD�K*�iB5K)���T%��D�wqy[~D�_�[I{���8�.�'ѣ���q�����i��W71�Њvb�V"j,�����_c�O*�xD�m '����2�V��wxS���Z&gn@��͂b�%�����`����3��'�6��}8K�@=���*R�`�}L��'/0�����%Rd,�0�Ŀ9	�-W9��|�L�1MF'��&,�w���~7�Bϯ�I�S�&!Ij������<�#ȶ�����lg,񞯐���|}/���8q:���2;]Ax/]��X�?�r��l��U-�at�'����Vɼ���id`���>h��y=�C
NnZ���'��.��6�Gy�	�n��؞�+�����M����J7�U;���n���2Y�ƾ^��}e���\0s�E�X�{ul�����n�D��D��>B=� g�e	�����z�>}�	�zy��J�����.$�3��^�F{�Hb��IC�4�1l��q9�͡W������mm���{9�|bXpD�[��l�T
_}�Τx������p2���ַ;pEz^��/9�dΈd��wr~Zz�)S���T����S=���k@g���%i{��#�$��+�M.�����{U��)T:ȶ�Z�	NYy��o3]8�0"�}��&:��y��쌇'���
i�μ�����;�����d�(#�:ax ��7����$R�<�Av�B��* �K���}�ݞ�{S�g�%)��(�w��/��S��˅����� ߈��O��A�B�T�I� m��{x_��q�B�؞�v�^��e�����uC;_��䕸5��y�t[�����Z��=���뙩��
�?��)�+���#Q��#���G-�@�;�mU< x���%t��^	�g��W����ޚ���P	�p#ɼ40����6&Y���g�����p���t3��~�e���)Df!쨳�l��:CCݫط���v�l��q���Y�'��*ԨCb��Qs��]�#R�����,�AJy�C㲆 0���'����ο�+Lė+MR8���	�:�(�E��!��9h�JL��^��{��d��<�_DU�X*Ț�hM-�x��m-3e����C�E��O�.cn�m���,7�3���\�:�QqP����p�L�%��	����"�}L�w���ږ����]F������R�����~S:��Rv�LA�`�,��Wjd���r��.MO�Z�KK{g�t�S�$?�� :���b z:���1�o�XU�`���fE2�������&"��d�	#G�6��-T��Zj�M�*>�C�Nˬ<.����?TxcP�&�_�E8��tu�R��1�P�ܜ"���s�Y����d��e�%����� �,²HÜɰo2�ü��������-���=]@��0�fTra�Ѡ�g�����]:�������\��9�O�Hg�ᑥ8l�2����}@�U
�P5��-����D����|�Ҧ�O�S���e�T��9ql�-�b�����y�#�N/7���\�=�*��{��A�AH�}����2!K���-�4p&�,�؋M_e�Aˍ|G|�ĤPтS��oQ=/��I�!��r.U��o�@
�3�W�&
����2K����!�""��L�C'��xz�Y��u�L�� ��N₏�:<�Mí����O��	���/�n�?��W�_b6������o ����-l~A٢Z��Փ0�cU�,�G3f+�Ov��ʔɥ��P:I&D�
v�������.�_���i^Dz�)3�W*b�w��/��>nKo��:]M���65`��r۩]���G|��G���ٴҴ��X4�+�$c��7�5D-�� ���r0ܬ~'���fT��c��&$��nR>����q�)I��}Mc�I4��԰ʇƢ�)���yU����|�y�(�/^E	i<�G�t����[!��i�������2܌�P8����/,ļ�ʭӔ�q	� ��׵7���i�,�}�Ղ�dOuMsu�?z��^M,҄W;Vz�~W����:ξ��l�!�A@I�% V�TT�!�;]��Q��6�j`�:]^'�+À�v�Zp��c�M&OTsEw� �'�P�k�7�CM��ؖ�?��7�x�5(<}�A��1Ȍ���*pf$��+��^ޫ����Z�k�Ai�$U8b�����lU��D$p��9��|}�KͱX^���]�ld��m5��{<7��,j���Ł\���V%����;�F3Eġa��j�1]; rՁg"���0��|�E<]�-��AvtNq�u+�.; �W>�ߧ����QD�f�6�٭�f�2����Dc]y��X8���6<�O��?�$+�(����J��
��] #Ʈ�@�!(O��}�^�3��.��"�Pzk�͍~n���5�0VN����YT�Y�)ɋ���g1��2�:uMᛈ�Ff̪�"�]	��`<Ӷ���a�G�Q������K�2�Y->b�jA����ԣMI�"n�ؖ�3"+;����%Y_��Sn$�Y���c-yrV�[9�R�)��:������>�C��(;\�sfF��[$�7�Lw[`3<����;�+o�G5�߮�̓>��Ӓu�*a�����gǀ`�����r�;�k1��DY�����k᯦�r<��"������{x1�*�ḕ�"B�!H�R=�&I�T+����o���,�J�����,�N�F�6��  ��pnX_�6Gb�V���N-i]��?-�+���#20A@��m�q0���������X2GDV�<2���$�x��s��|��	�o�;@�!�,�Z�v���m��	���y
��Y1�D�C�gh$©V���Έ�V�X�E�"�5V?ʯ�x��vA�H����5�!��E�~!~�9��4d�&Rd[��d��P�E�i�߲f��2�,�q2�mJ�	�S���#����=�AM���~9��u YD�ԍ�VH;�˧�=�?Zs� ia���FO�!����F�#���i?I�^�,�m�RH7�j<��y��ި|����1غY��Y.͇��L��AӸ/sL�N�bY%�U��@ʬj��ڭ"fM&�~E��~��##�>K́y/�xc�Ҵ
+�
�~=����?M�z�L9�A�l��S�[A�pC�{o���=�".&��Y}�q�=5���~���'+o�uݴ�7��3���1�j#�T)N�-��:�K݃�uc:0������9�<������*���}�d��"h]F��C9����ނZ�IdE��Ĭ�jn(EUj��9�P��(����B.q�q���
,��N�]��3�]��F��" -ǘ5���Y��	'��{?�.-�<n@E�����M�A��&+��>���M]�#����/cY�*���P�8Q�%T ��	����nF$T�wC���=k6�?r����bl���U�I��ғ<~�$�,�N��q[�:跣x��m���oդ�-ґޖ�Ne�.nK�m�����>����v���o�&�$��n�f�@�*������2X��t�	��M��R�]&	w\�!���!*��CEc%�!�'�~�ua���������nS2�Io�E�c�����v�����ɳR� �0.��ċ���y�`�`��萫ep��A��J���z����HL.`"�샟ztdJ�� ["��jI���|�~���|�rΣ�w �\C)��~>P
|�	��Bh6Z�*�����?7$BT��_d��߄�,�c���$^�)r�q�q��x�t�ʛ-XX����0=fLH����`P�kod�}�Az^���DH�ԓ4�6;fz����-�L��ۋ���H4:ܙ��zǕ� ;�@)�~i���N�Ls&%�i���<欽�����N�d�O����B�t�[�dQj��$�bRش���%�¶1��ju]<�����ȍ��C�a���T������*{���<�W��8 �UB��r9�� �*����Q <���l�9����ɸ�Wo��#��W�6ޤt�@����W������/ƃ�(.'y"`�@I�����F��fv2~b���e��@�* '-uT����B�P�&��4��\U�sL	�Y�fy.EL�;�Wd�-N����(�=�f�I@�@���,P˘EBQ�]��*�5/��̂T��m=��J�'�o6f�LWA��Ql��tב)~��_%�C������M]"�%`Pݜ�`;{L�a��@��Xi�}^��� dȯ�猘�2|��xaO��-�ų�M����UM�:�$`��SZs~�J��!9���
�Hs�o��}U�I���G�k��ї� ���4o�^�y��y�q*�L�K����ڰ�>��w���\��?���+�sd����I�+d�b #�\R?^y�����: ���ףhp�ROi��i��옛[�3��!�0 ;�\q���c��Fz�����s'޾�;���`|S�k[̓/�1n/|���/����ވ��8�f`��6�CyH�5J�N�.h{ͮ�{m�4Y�!XOK�eh�H�ъ6>�Y](�U�bύ
B5W�F��Q-��fD�$��\�}�+Em&X��},��jM���|��B݉�+Vz��?�e���;�s��/��/�
��3�ժ$'���f (TV�94O���J��G�o/VW|ڌ�x�[?vi��j%T�r',��)Y"_a	7VE ކ:>M��jtr�8�%���N_�N���
D����Ú��F�|��&��'�ath$�L%?�A��0T<Ӕ��P��r��<J8�}��h����ȹ�"ʸ�V�I�@��?�:͡�
r��H�"x./�^!X��r�E�����/�FEY��i[6��~�LHW�
�gU��kqy��q�/�'/K�mЖ��[7���=�Y��R�d^���I�k�W�^�NA�B�2�`}�1h�AI�p������A麋���
g�h)��� ;+T rF���
=L�2J0L^�c[���x���r��C�k�s�t&'Q!Rۣ�::��/6l0�P�(K�^��U�$�2������k��Q�G!�L���W�x�l��v�۾����H;��������'z�}� ��A��:Y�V��k`�Jjp���A��r��O�A�7
p��Ͻ��y��������&��i)����]��	�&ҵ�~Eߛ��8���mNhR��_w�8�����[Lͳ�o̸8��4ܳ���G�Ϋx��\=�����V���'ٴ�a� |꾒I"�pj�j���K8)w�-em
�N~��K��$�R^P�4�)tt��4HD"�A�,��=���� �Uh�534\���XaZ�S{[�2?բ=Ei���A�2v2�#�rq�۵x�����*�!h8j;�o8.knܖuE�z��ޏ��^�w���*Ƶ
�����Ms��9	י��a�Nu�ᬪH���pe`�Ǘc��-uVs-pxI8��'�'{��R���������g�ط�%u_���]�(V�s�1(w�����WKn����yt�,�$��Ԩ�%D3�P8ba�O�N1L����lԃCC��,L���A�5�ؐÉ�Sb��8�fHI8:Ȼ�\M�TS�K�Q��+���c��*��0�����Nّ�q�ӄ-#�]1��q��J�<�hQ51���?�:�T%I�"����9����¾*Z�\Gpi3�d���~t������Hl�0�J���q~�{�pnP w0μ&��!��S"O2�Ukg������m� ��pnJ�ݖk0[�K��cc�\�s�y*>I�Dv��a�+-�w��㓰��:.�#%�kͬpO(�$�S��śQq��P�,���R��l�,TK���b����&g�r�Pd��vLTx:M��f�zqUjP~��[R9�8�-7ɞŚ�&�����w ���0�~h�I��q:M�@JDa����c��b�O�
{�$��ڐ��]^Z��h���$�֗�Ѽ����]*߀+�l�mB���ꌔ�lW��#@���~�\JG�^\�2��0��m�S�m5�P�:x/�M����I���ǽ�Nl��lq�K�� (f~֛����R�m:9��o#X�o8�^yD�wJL����IW��/��ٻ��
R�?F�^��[̢���=�z�R�h�����Z<�̿�T&Ld��Ll�?��B=W%T�%�.>���滲�ə��/��Z^�;�Qr8�i��t�w�-��~�{��Hܖ*�q(���bx�ǵs�i�o�> ��/cyW;+�eG�S��Э�eiB\����+�դ??F���wn�[J���.���hR���`�%�����o�4O@��nw�ľ���/뫖v;�q��[���=vn���	m�S�(�C����l��@#(=Q �f�1s���%	�M0JZ>5���D�H�-��1��{���4���&�h�6��I��G���r��:-z�bݡ�<&��F�
��^U�����1S
��R��w���p�Pz��5�zGh�1~J�n����_��֏bO?��%���q�[��&�^�nW�z�X�:�PI��u-*%b�a��������IҒ\����:��˓���!�K� =a��_A�C���k�P2uU����Q�甮�(�Zwu8��i8##���Y��8���p/�7h��lb9h�>�H}�T��-�L]~Qx��H��i�C��^C�����*���avɤ�ԀwT�uTB)hũ0� ����C�N���������&�m����aaz�̰֞�u8�w�?�,�eLo4y���w�F�1R���=IY���1�KN�:ɕ�U�#s��7D�,GT�h9Α3�5W���� "W�!�������{O��J��yZ�򳩬���X��Eo�龥�f�"V����ioq�?�J�^#����L��N�"��и��?7����'�߻6rjZ����yȻ��6n�C�8��͓vgW4zg�O����7����=z[��n/�����&��sp��֊+�ۃ4y�&�B7x���繾��et��l<��F٘�T�|ɇy��5��v�0�-�P,x';�q�l��A�h�	��l[e2��l�� ��ۛ�+%3Ű��3��Y���G�?��סcB�k�X�Ѧu.o��b���X�o�Q���sa�aև�Q]%;�&R8՟C�c�	#"W>8�/��~씃nfg9�) 2C�N�k��(��)�U| ��Z�Za�d��r�oj!�M^x�X�
�yh�Eɑ�Tȁi�s�n�(C/'
�$�i旱�s+��|S3���9l'#��o��y3D��Q�ܝl5DQs�$���H�x8��)1��h�(���t�%GlH�鐠-h�q�ly&������Q�tr�Lˡ�0%>����H�6������WO�"��e�A�8�	�׷�b�+<'alC�|��`;F����e��e�(�Z��0T�����e6-�ӺgW��q[v��=�'�R���@�4�V٬[���`)Fa�Ɣf��`�!�RW.ߖ�d2��AՁ��r
���Aӡ��<b�W]n�����͕��=�1����/8�er�į�:��)Ӆ�r���nڒqp�� �N]kX��UQ��*��Mx���^_&u���D���8���V����;��c��g�<�$q^C�wAħ1~��R��!�#7�W�,u��q�$}��i���6�5�u���+×X`Męw�>B�[����V7H�1-�z(��G⯶�3���m�|�r7Ƅ����t��>&�F2G��g2�¤#x���P?�0��("�UH2X����|X�G��%�Jy� f]`]0����Őo#��&.�fc��B��gG����nD5O���z­T$Z��sw��*
�b��P@�Utz)���	���o����z��ۍ$�G���0�Ȥr���Q�%��1
F����Ķֳ�3f���=e�Vq�����I�]�v�Ʉ��[!�p]�M.�Y�%Be�� _��'8��z?9���Iq�D^P�[T��2ǵ���!%q��0�׆�aq,��@���kq��ڥin�/�T؛x��qF�G�����yO.Q��� ����r�F)-��v��,�k�8Ю�:>B�R-������0�cW�+���CRp�Ufg��)ܹ^*�y��گ46P�������-g��E�$-�9�Y�I��/��j����Y��>�#s��OHԚC<�;��Ph��U�|�B��B�ͥ����~Y�l7Z����[�h����1*04�Ve�Uo�BH�|7/��������M���Q	9U��JI�=�U8�i���B��ĸʗȘ?q�8�r�}-�7�׀sg�
�����N���15�������I��m��^�'�Y���aFE��dSU����✐�>������c�����)ȑI�����t�@q�w�/�x���@�r>�T�$`1FVJJ.:����X逐�"&Dm"�5}�D�J�XJ(_�:S����-�YQ�&t�-H@0u��ɹ�x�PT0+53���桘�g�?v�P�CQu�q)����f�d��Nې�����s����`OO�U>�bX��ج^�a��ʡ�������ID���K�Մ*HP!��+��nD:�����Ѯ8� �t/h)a	��Fx/!8J����E�c�!�;�S�T2��bE�g5�o&7�)�m��1�zd.5D�_����r,�<���w������A&��v���\�n��W���ʠ�p{�h�d�Q��I�G�&s�0���Ma�5H8�Y՛A�iO�7����Ih@d&��.ֱ���YBD�-18|Wg�Y��-P��ç��Mw��J����(}�,v-���r�M �b��P&�J/�)Ϡ����
Yl�V�0���V��:��"K3T�#�մ��Q��R
����'�DN�JGA��0�6��5X]4�G������$!���Mи�ww:|��\w�אýp�-ӛ�[E�r�k(�Ջ���jU�匍�).z���B$9�I�~6Y< �*����mi���M�����wK��Ы	W��}&<��W���\"X�}-��>���E��&b�Y3���w�WYb�j��7ᯌ!L�q@%(�7���p�����c~.�GM-x���y�������XRE�y`�H���	Ȓ�mH�#�Oz!�$�4����;B>�f;�h?4����X$��0q�#�pvq^��@�},���� �#۝U����$|�លv���-�4�ᜬ���'_%��R�,j�V7L���̄��\�A<j��tS2�u��h�j�?Ɨ`M��Fb]f}f�t+$�8aj�uAҋ"�Y~��Ky��/#lIƿ�2Hݎ'�H����\o����]0ڟ@�|�C�A�O�Av���O�/�#X�'dhN���X흓�¼����@���-�f%��d�������zM0}����W��͟�䘏�ת2�>}	��h�HU%ĿR���|Ag{�$,Jz��]?k�:�-�B#����B1�bw�܅3c�PF�ψ��1:},�O}2�u�+��I=}�dBۓ`K�Ƶ�w�콈S�3JD��B�h>�$zo�Lk�@�]�?a�wB&_��JE�$��<�߅L����Ze���%�g8��0 �X��ԁ?R��/�HC=E���	� >t�$n��C�6yb�Hm�/�0h�p�p�c;o?C��"�z{�JI�׻�9�Y@h��u�5 6h&X�lU�詊Eŉ"y�d�M�ru��O���	!�[1��z�`��D����v��TU�Eyq��T���?�(���d��x�K9�2���M��j4�O�{�t\��{o	Y��}r�>����-->��iC�S8FW��'|Y8Y�$��c�~�e��]�x�"��}�=p�J�����3��7��"]��������Yє9����2I�k�;��&�E��r���T�;�VLg�a��~�'DHW.�
�ή�!�����!�1�=I���@�uI9>�}�\�4w�N�ԑI�j2i,2P�z�q�޺*�>�r�XR�����B���F.�em��	瀁v@gp����`��Z���)�fY��]!`A�@+��	�k�p�ࠋ�"�Wq/w�HJ\�#�V��l`֗��5���5�D4S�*�w'{޳��WifV� 7�L�liFnU�5��CK�x)��u�r6�$�k�Y��]
�
������ծ�#|��>� rQ���EAq���U����������X�Oӧlj��,d#��{B�C��o��I楰����x�^Hg�M��ᅩ��8�vӾ���͸��@����_�qg)�a�da��z�4�_J�[;M����+��Z*LJǼ�ɹ�=G����V�J�v��4Ұ�;Y�*��'E����X�%�8�#���[�u�}3�%o��<�t�_�O�η�(��C�}`Q�`'��79P������C����!!D54�J��.�Sv	y�1~�_��\��[���W�(��jS�@�}u���ޖ��nڥ�;�f]�V�1+=�˛�ph�W��P�wH!����g*�'�sJ 	�TנO��>D�X�]o�-�Cb�������<�}o���t��y|�~Jt��+Z$�\�B�*r�����䈷��2Q	ɅI|��b��pqN�KiX�rp/�N?�,��M�,�;�8�.X�?�(���ᾮ�̖ctS��1�fA�I9��~�͢˓LSy�#zћٹ���:�]'M�ت0��c<wW�G�14�'DVe���.zY/�w�=[�d�ă��0�����&ƴ,tE�&)�-yZds�"��O��FT4�:F�khx��G)�<���N�;�����M�Y��8S���X�$J�t��m!&y�CcJ�v?����T�oJ���'����O�e{�W�*rOe�m���	��Z�0����a�����c��ڙ
b
�9r	c���Q?�A�O<\?e-o�Atp�ܽ�|�c����\�x�X�Ԯ�q{\խ�b�E�:RЬ.�D%'����6b�QG�k�vT �fm�18�������-=t<G�g�ά�!��d#�_�V��I�`���QMbu�0������m�V���ID(>�|��?$Bh�ϫ-T�3�8��*�
W�=���h���f1�?��i
��?.y���T36�6�ڗ�Ah�r�Db���ľ����*�Ij�������$!t�ѫ��eC����*�0A�.\g9�΋�t03�������B����3W���{NY{�*I>�}��j��	Y02����X,]P��<���?�0�E��jH�c�W,��,'�.��3�� �ʹ��0!B�W�W�>�Hz�ZK�`��S/G-p�Z�F#��"�w�K:��V&)\3f�]����Ngah��| a�W��6���;n����UOb �D���/����*ݠ�0#:Q!���,�'Fɟ�}�xR���� �������1@���02:W����k��b�x$�l��sk��[Q���'} ( [~_QJ�JMs�&���� ��q�]<83�f�����|��(l]6�����`�}���^�tz6z��Onj)Q@f�}B�!$��쳭���(�쾺El��!Q��d�֮{��X��u*��/� tCt6�=���r�B��T�q��/�ljOu���f�T��4K ��g��:l3M�6�Y6!(������N�)�_�0�s�_m'/D)n����IUu���,��������a�/PQh������ɡ$��0I�dQ���c�
�m)_��S��F��7�V�"��k��Ͳ�#p,k��`�S�/9�%%�ޒ�t�ꒅT��������g��hC�Z[G�Px�^}3��˫��N J��zn����NQ�r+&{�W�,��U.e���RčkB���������{��.9a�Ϛ�Y��)E�4��5(��JN�*fl[S�h�|*Ѷ�T�|��AU�#]�c+����0_�Ym�DJtԼ�E�3�CsSo��G>�,:�m��X����V��1~kgޅ*7�W�y�.�����_���b��cɔ�(Q'�,O��xneIx2��|Km�~��9���Z��NlW��JTW��I�0� �y�$��J���,�����9�XW�X��'�K��3[���Tg{���["�]S�~���9��Ƒf��+=9���Z�#C?���X�#ͻ����=\߃�^����=OO�����w��Hʐ9A*�8="`'�ZT����ܑ!�E*�>t��sq�a�U�x�Z�/�D}���^���	uZ��j�2x%P� ��������D�p���b�4�ƼA�08.��M�i�y�漋nTkը+DIA^C��Y�6�W�5"V,Lτ�j�	0���OUL����h�s���j��������r������Bt��P:,��wT���x<T���>�yT�y�������" +�GOj#��\:�wq�m����EVz��1�	��A9�%�F��J�릹CQ��]u�A� �(�VDu�7F���y��)�[P!:����R�Rb�@��5qVqz9mv��?�o�z6b���mK`�d�EȱT�tK����2QU�c2���S��oΙ���ծ��,�sT� ��Ù�#�"�wT����pZ�^��,��J��r�`S�j!igJ����~��9�B����$-nz���wzd�*x6���eC��z�f*_"���M{[��1�}��e��L>^T̽��	`�\O<#Н0�E$1�"�[��rur�X��'v5�H��q��o28�I�gt+��]�QV�ISy^�7V��7�]��t�ႍ��~�w�Aؖy�������3�԰��Pm^#�4N QM��2�ǤW)��1���@t6w~���(�����*=AJ �bխ��'�2C��UNϞ�*�P�Cp!w�f�����e���v(��](L(�(�tc�_����X��Z�����B�J'�����潧�T2�d3f��We�4����HB�XR%8�¢�W���Bm��2���]��Bz�،��-v4L�����Fumg�g���y��B�ݨ7�cY����!��R�'~O/��C�������|_����X�8OA�g��3�w,P���/�3+p�(''<�O�&Rm2/��g��F�g��Oa�
 7���+��b�������U&pz��E�G���� ���S�cxM��ޢ�pC+_R$`���Ž��f���vp��Ja��0R��˺\(�,2г�у@��zyJo�Z��_��^|�ӭM���A�1*��4�phh�M� B��U~8�_�]���9�":�e���Xq2{�Ě�l�������vH2�������.�j*g��~ٝ�p3\e��s�v�9��╻�A�~���Zl;���%:N�H�k��8X����݅}X�6������%�*���>y�}��5{ +�Tߙ��1�+^�rT�G�GJ��o)�����y��+fYݘ��^6����0l��5i!�sy�M��V �޴���:s-	d|B}��89�P���C�<<�`�p�~ͷ�DEU������vu�=�����|���V�H�c��MHڨ���5Z�:xM��ZL:�u$X��$�l��	?�A#u��r�Q��G���0Mz�|X��@�;F	*��!j��M]�0R������N^���/)a�0_�HC����>�7W����S(����VE�����{|��b�vE���ڸR��զ��8����,�I���xLA�Bى���b��z��F�q�_[�es�#s��~�)�H������,��D2�c�7%	�u��4t�/����얱��;nS�J��v����Xl�WhW��W�7�wy���l�<�������psybYK�O ט3�׊Z�ڨNJV��|�H|���"�����j�Es�v����!;��(���!!^,Fgv^����b|V���ؠ��	Djo`�^��և��L��:
���wtX9qc@�����������9�0��� �@�C6#E�}��Ai~�>܄t�����ͱ��9Sm3��/��2ȝdT
����E{<�G"֕���r�I��+0�f���G䴏������?;�I������)5.� �0�(�opLP�񽝑%w"wv�c����$��C�;q�a��ΕE�iTi)��,
??R�b���:��U�~�;z������5���xU?ѷ���l|�&u������Fy�0 tB3�i���ώ9��0�F�hD��l���(��y����Z�B�B��>��O`���:���/�"䮤�2$I~��KNc{ԯ�XD�E��ݛ��3�0����CS�1�y�=�߰|~Ⳝ��A}+8��0��D����2�ד��*��ȟ�f��'�5�2Qҹ��o�.�ca� #��Q�c������=���lfH�6��7�t9ڧ���q[;��*�6�GDZ��TO�χF/1㧽6 ��n�8g�!���d��F�D�@���6J�5[��Ua4�
�yā#�8��Mt�UKT�%K��o�<�f�,%/ߒ��v��ww�c���BË�Q ��.�{����wf>\��	�;�t �����5Y�Ә��x�ک �]C@�����ōEG� m��A)SA��j9J�<8c�,6Ĵ����L����"���\��A���5|���_��T�z�gx�[S�e�6�t'�\��K�~��QSV^h�Zn�=)G��g�X�WW�[x���>�KW��1$����Q>&:iD����.���ȏ�"K0�ȓXQ�������8�gg,�#c�|�"���κ-aEOY�����y����$O�d�c���GV{,{����Eb#v�7�����&���)�K�sv::�(JS��{�����Q�[j]ξ�������{$<n� G�čѪ��C�λ虄���1R1\�r�o�PU��A�	�����)ʡ<@�k�������o*1硍O��0S.���ݛ�/�S\�>��=�s,�P�8_�JcN��l
��\�wݘF���ԋR�h�	��b�O��]+U-HD������*�~a��4 M�,@{Y��`��� x{��݂̒CT��Ҥ��εu�ᘩ��F��F~m��1�^�ݠS��-Gck��sV��h���ݞ캕[,/o�l�B�zp)���_GL���l2�SZ���Q<��;-:�A�\���7���Ů(��؏ӷ����������D�ݧ}�E��#kL�����O�Z3��Ϸ��.�wB��M⮠!0E{#���;���9��jꉙe���뭈N)P�-�w��'�����tn7)��O�D5�;J���E��fD��(�⅜��?�0���.��M��Q����f}~ʬ�A0�K��N�>�f��\�2��{iǩ:Nڗ^��ɵg���o���(LǨp#�"�g&� g	��=�K��c�
2I���pd z��.,~	��'	�� :m��b�J�$�XI����}�Y3m��(��7t4a���}sA��fs���`j���ۓ��4o��[�;�Jr�!��lwi)���|��_P�5����"5��[�����,�&�/��,a-Wh ��ht��Y�ӯ�E.�\����a�H4�e+��s��-`���K�{j�5��)pJӽ�����'�{���˞W��Ww͓��=G�%�X�h*e���`���f��u��>�s
���7�@��Z�=F�YPYJF���x�]�C.�3�
��GYb?��V!�S�i���u����v�YF���+���:k�0Ca��+XL�95v<�"SRu����ಥF�I
��C���0Ȓ�ő�6���|��\��QDik쓌�r"�b&v}u��T�̂��l�!%h�m�)��}�*�&��T���Gp�A)L]���L��(s�>�('0ӸvAf���Xy�a�'��[<<�b��s,m��E�ܑ
N�Q�T�� ��bqBx��jw�ٵ�T��T�.�2�-��vUkV\q>�9��#����B��5�P��}�My�H��a*��$6`�<�U�����H�=��f?f�`F��{�G��aZC��F��~E�r��[��`1�:�X�$ɣǽ��S�RU�ɢ.#��~��y��#�q�i�һVG��p�ό��%K;�ɔ�[��|fo���s��etzK��?��JŪ#�'Q`m��sIEB�sHL��O�sb�J�RG)��ppiӨ>�)ڲmE3ĪD�2&c�}4W[
����h|���LP@tw�����=UUG]`�Jp���n�ឡF)��WG�[j\�Cҙ�?:^�o���Z� ~�8W����� �|���>+�Ng��t���F ���_�
�����Ê!�U�M)�J�.ײK|�
�{���z��@aF�W���9��H
�ϩvt��a��_�>iT��K�e��CP�hT,c�i�^��D��Vj茀ձ�G��w�ȩq����a�b�I��q,�Ӡ���
,��}�De�%�Jqb��|�6��K���b�M�_-5+��4ﺽ;��v��~���p��gj]���ɑ�	�K3F	��*I���"�ڬQ8ݹ{���Mh@*~.��:R���K�r&�.a�[����@���z?y�x���Jj9b��%�9@b��S��O��xS�<��(��ټ�.]]Bh����8;d�G5'3���fW>�:Z�[nO���fՒ@A����/��34`���3d�J)��Է|]$�FMJ���9�76<wjD�ua�K$B�����L��q\��Ӛڟ�A�׽\o}O�
H�7R�J�̗�bKR|+��=���>���ʶ����zp9�9Qa-�oK�3�#li~;dJ�_ǚS{D�Uh%ɷ�5��������t0��-�����t��RFu�[�d�{0���W+��#�Ri�;�F���v[�X!w�z�jt���@E�闁��g�U�a�#�sؘ6��z��)���b��S��=��ǣZ��s��H��c�[���e�E�PY�К�O��nM��n:w�m�M���MŁ;}��:��k�v��l
������ba�}F/�`�ؖRŅ�Cy	������s£m~���?
��ɫ6����p�$��q�Zn1�Vi�����J-��C�@�g*FEG'�V���T�BA]����h	қ?�~r+���o�������9Aq����5?K��l��Go$䭘��?Rۅ����;�Z! �Z����~��UQ"����M�~�y��Hpٟ�xL N-�b`��'�cU��%�)Bآ��[���3֑�� _;�;w�<�pMo��+E��2q�mo�X��|�<��u�b��w�!�VT���b\���{Z(�kT�b^�| =�����mӇ�� i�����F�Ҟ})��:Ɉ33��`��n L:�k$©�	��#���i}fM�5���"��+D��єݙT ������е�@O2��������QvN������wD� �<���NB#M0Sp��˪��¦c?&�!���OŐ�>v�Ĕv퀝t�[
���J�^a��k��G�P=��F��$҂�
@���)���R��Sbnp��}j����̍s�̿-	�����V��_���Ǔ<�k�,lds�� 7m��f�B���G9�JsB��:QYn��+�i�aт���4�(���;��eV {�wt��^*��D�_#��������2Ƽ~IY�^<!��k4�{���F�����yQp�����?��lq������2���@�I?D�p%�WŌ_:�~E(�w�~mU��4���t��fɓ�?\��暊�iR�Y�W��T*q���T�S���A{5���4���)�I<"q�FAw�o�%݈ưwp*,��4�o\�]߅��H�yZq�c�����y���7�Z�_�s��H����pu����=��	�2(h��-���y�)Ĥ��M���
�ղ5}�&�����t��l+*�O�T��[�c��\��Ix�,��#Q�;�ZJ���.���M���d0�@�R��ˑ4ɉӠ]/�%�V*��u��[]HP5.�D:��d����g����p���'�5��!�(#���ؗ��Xq�{�$j������l��U��&
ѻy�2A��(�%c���U�AS�Y�Zm���D��1?y��f���ʪ)��q�ϳ���ʜ%���5�,�j-fR*�}�s�C��!�o�y�k#���|�Kn]�� ���ȓ��$� �����d�4óƠ\�ރ[%ćv���
�7|�'e�lU�H�+��S+޴m��GA������N�[��X�;�Oƽ���v����� ���LR��{1$5�aY�Y�z�UUG�؁�᳎w�+QV���T����gR�0��nK�{�Л�q	��%j-����2ͤC���nڄ��v�u�����nA�%��˱���oԤ�6eU��J�T�o���Be'���_ƻ�V��9�V��=v��`d�,N�é���i��|��m��W�L4��֖.��X.nJjo<6����FӔ=��C~1L(0����1���&W�I([.���OxQ7�/�{::�^�A�e���Fn u&���\�jC��{��م��*]��@`�3F��c ��uȑj�l-�!,��}�ȹ��@������N�PR�A��-�|����cPQ�:�\pB��������ȋ�D�i*�:�JL�9�3�� ��5���s7�H ,╖u���f���!��ofQ'�R�9���%��yܐ��G�5VTލ�+lD��9�>Esz�����N�%ұ�>3������ L��CsU��U����ط�~3���_�5�Y�N��"d'��1�p*��l��w�E��_6m(+Ѫb�3=]���VMJ�V]�N@�g
X��J/'u����)�<�{ ����O�/��iWƳ&+���q�����t|dG�N��w��2zקF��tZk�Tfp��˻r��_X������U�ig�)+y=����#(���W~�WŪM�29�Y��uD�==�s�K
g�,�"����� ����aQ�Jx����zYOb��]��Ǧ��*~$��"��1����Y�2�M���ɇcS���M��Hn ���E��̭��}<��O�鳞:�#�	G|��ƐNV'`��0��u,�m~��@��&�4�2� T2J�2kCE2��F5Ð������EA@(�{䣰'�E�\2Jd��R�Z�'�Q,I��A�^�#�ǧP�g���D~�\i�]���G�B���|~z����y�A�,sQM�|�*��0�[C_tg��R2n|�[1�EB�� �oڽ���|A��ŗ.v{(�0��lsw=%�#�Z�Lkk���~��IT'Znߘ��{nS��4�a�30�ϥ��+U��E�f�	x�k�D^��\r�R2i�(����T:�W�!���{�칠����r�$�2X�%�����2�:����7w3MJ#I��e����ˡ�6	]��(wa�����>�����K���+�+C����~C~������E-�t��.��r5��cy�z]2�9��^��T�$=z,'�p��yd!�)���Q)���7�L�
��3�{Q�)�8j�ɞ��S����s���B3���a��-�%��D��=)�?a�B�e �:�FZ�,��KL�wCɌ5�^Rۋ~F
��4 �{�Gׯ-�9=!���%S�k�̍��[}��|8���u6���.<g�|�{���GR�y� E�{E�.�ӞrK�Ƹ��60��6y,Pn�{�/ԩ�5��˅>(������jl?��9֟#�è�z���O�P���"JI��Ǟ��|�"G��0omgg����5�HC�;�y�]8�$7U�-��(:�(�P��W���N�ֵCMpW�1ҕ�m�Gy��9���jrU�(�e|��i�ف��r�����9#"��$s�b���	�h��1S��x\�B�f�|L!�U����y�>�&d���V}��Q�Z�N�9���?��v�MkG
���L+�D���v`�ǲ�R.^�2�ag����k��ݢ��b�eI�����l�������̕X�EiF�G�E���?u��n�E��7��ϊP]�4 D��y�31�Mz�P0��9U��/��8����=��\���0ZE�?f�	ü>$�|�-�R�@���=�Wz�-�kmM�܊{_ntyo�7퍽{� �`Do�F�����Ds�ZT��=*�X ���S��j+�������o`w��'���>pOc;<C�K���j�g������8��_��$���Ef+�q��אhcP�P��/o7$!;*׋PjN��|�n�qx���BZRh2Z�c��k����Q�<����l��'F��h@��#)��g�?I?R�l�{��#_jVS����)i�z�:ܛ�G����^b����D�a"r�鴦�8U��DB�m��#��ge��ϲ4�g96]ϡS�7�F�O	��H�]EA� 9(�\��Ӄ͵7���b\B�,��_]�͗�@�٩O�{�4E�ۊD���F'���?a���,jf������ ���%�[ӋP�n��`0��d�_4{F��f ��&e��)����d�^!M85������u�f��3�{nGgrj��R�B&���g��C�A���K�	~86�E�gL�j�IÁo�A��ޕ�:&�x�����x�Tz�&X�R�T��U>��.���8��,O��ԷUd^�����������EN�Z��A�l\�`��ݿ��q�h�1�,&�f�b��RYY���$+T{��T$��B�VaBă~�#���O}{H2.ݤB��3����Q禅 {_w,_i�����4i�E;H�Y����:;ͱ�����[�np�3*D?�6�F7����>�uw��7i76dt�T���v�';PU��?��Ϫ2���.��Ҋc������:W�Y��͓@*^X���/w�i�8L}4YC2�+�I<�u]�A��AM�����<�}�&=�0gh�/��Z�~f�DM<Ϣ[8�MIK�*�PE��
��p��®��-�6߼��}�\-�$h����*��{e�O�$�#�g���yK`�H��U�9Xf@vXqɊ{{4�"�s4� �v�m!W&?[��	���r@�$_��%х�y5�^��2[0�pB�3;��������m?胗,�m��o�����p��  O f�j}]vy]�$���\�c�PM������ ��D#�?ÊZ�n���qrC�_u���>�Z����J�)�u�wF�t ��#�	'uj�2��.��XJ��%`�QA�k�(����9�u��c�nR\-?]�=���DN�C���\;�2��KsQz�g�+}��Fm�Ï���xܳ���6Bx�w�0*L5�"��iT�f���A��գo$���7�&^����q���[�y�`�y��֟��#-�H^m��(�I_jO��Es��
LL�l�f��;�e/̹�rˠkD|[LwKC��p�e2�zW�?���o'�j�#j����R{�(�e�7g<����&zq�JA�V�A-i������J���f9Uo�E.r��9|mC��o��b+ɺ�K4�Vs�smG�]8�pY��k�Jm���Phu�p:���<甃��(�ZVq0>��k�Cl����%I�߁CtR�z ^Fj�O6ޫ��?G�~���4ʉ6m՚���eo3<�lRd�xC �Ѫ�|.0��>?�X�k�N8�Wjb��2Ж{%@Ɔ��|7���>sW����p����UH�-M!n������8j��L�s0� �j�Y@H��L龣X����e���h�#�U�b`i�����]
.�}���0C8�
r����%��aUo����A:K8�d;YN��k7�')_Mi��>�Kl���s�鰋�W4'B����+�����r ��4���R���T"���|9Q�;ߢ߳��tp���[��"'�' �'�:�]���޸�r�R���O1��t?�۹�9�׿i�hO��L�m����-��C�F�JU���*�K��aC�(*�[�
 �b�L�}~t�ω�܂��%�!\��N�%ƣ�c�m���h(�i���Z�u(j��hb$��\����)�8�:*��:Y�/ȷ?�&�UdDELQ�.,�TJ�@�A�ȣ��� ��_-JnP�Yw7��Κ��4t�eQ^%[
��z]�ʢ ���md�%��h�	|:�M�l$��,����0�~�A<��=Q%�.���nCvS�Q��Ϟ�s�챌̉�6��+�����^3�ځdf�������=I�l���t�:�HFt��j�}.P�|�A�p��J�zB�0��G/W���[�1���~]�qb����~i^�;��3ua�%8����"��ǩir
�ۼ���>��.�����Ψ�`�*�fmM���2}`R�������Yo0pٰ��k/<�O��-�>s��r�C�yB�x o��6[t֋7���׺�Z-�;��7��y	��(4Cxdg��1�n,3cs�g���b)7�%�q�y�^P�5�]�=���j��^�\�5��&C�9��� n�e����)sWAR$��@��{�Γ|FA>���YU��h�.���x����t
�Uv�@yD��Ʋg��Ad���r��`��B���^�z�����à<~��
�=�b*��ow�������ed@�6"}C��#rKl-_F�.1�1�?��������19�K��v���277I��g�C0v�;�/ˌ�a[�Օ$%��5���`���j��L�}E/��HE���J�����֣�0`�zbdA�F/_ZB����;**������}�}-(��L)A�@���G�L� �	pj��'w��@Y{�s02P�P�;NI��Q��w���4�s}4�q�dI��r�V!��OqQ5��܎��U�����}b�l_v�`�h������m����aR�b�m��r��)Av60�#��{�o���}�0<���sy�!���}���&�v!�O�{}��^�I��N_r��W\m]W�MMY?������ ]�6.�4��kNՃ�H�� e���
��b�d R�q�2�S�B�s���ߢ�֗P��ݐ뤜�c	Q�,ύ���������|J�^�[�c?��&��y���|���\�]�Y}����E~��J��Ac�����l��&����J��&��������������nS�Vv+q�W��](҉�C'�3��j ��F�!����ܐ����ntD�+"l�ӽv�s�m��^"�z�=F#uj�Xi��po0�aiр(�f�������i�_>ϧe�*�Ȧ%[���|S��H��*���h��Q�o�T��;$ IY���i�)�b�۰�S�e=�BT�;���m�#+`>B�m K�Wm�AV=q-l�t7�T&2�C�2v���Y�s�58,�(��GR�[��8���0�%X!?�I�C=Ұ; �S{3�5�ǣ,%I�	gG��u?�j�z��"�G�Oq�M���r���J���t"����P�1�/)(\�D����Y�J����پjoA�9E@Wnq���qi�`K0���e�ب�?dd��{��� vF�V��։6����8�u��?���� u(AЂ蝵��CW�xZ{�,Ѻ��灅(�5	%�
�
9���K
3*���%QY�܄3����@'��3��֠v���x�yeEM�繆 ���rx^	����� �;T�޲.�F�T!���P|��˨�E��F�Zw��?���:c�
Π�T����E���#��'�}���H�����w���/�P��k,�k�#�I�	�����ZۢڃS���"��v�����XWJ,��f�|r��̸�1�a�c��MJ�������N����5n���@w�,;Q���#�Vw�� ���H7���kJ��\���i��=̵�����LB
��i����������'@��,�=��֓�������9� W�I����H����c�FH�@�G����Z��|�u�Bw��UP9E�I���
�}������$ ����=+/���SΩ�z��0�������B؁�Gju1�Q{�#���v j�|���m-��!
2����;�*X��.�Ri-�o��)�
��j�#0�q>�L��I���������%Tj-(��(���&�-������t"��wfdA��A�k��l!�b����[���R6�.f������9h��S��A'R�{�OJ�-˘0�tK�mfǻ�.�:������q'c4��4>�SR�S�[�6�Z4�X$����&��}�XT�i���e!)=��-��H^�<�����>ƭ��ki��.��ږCe���z��2k:���-ZPF�P��tC��`�����D��y�t������?_�.3Q�YK5$�����'z��>�W��V�$���G*�/
��uù��0Sx΅RMp�9`A��@�ɤ���aY*��t��mw�gR�x왇�S�+�aŮ̀g��I�˔jw�,=5�0����l��L��3pՀ��T��
���Yƽz~����w$*�u��j�91�1��T���2U��M.]n���<����o��x�^x�>�2?9�x���2�yu�k�k�I����j�Bk.�DR�TP������� w��U�Ӎ@�ID���.��y�x�6�N鬝��,��2`������XW�0o��۵/V�#���a=՛b�!��t�j/��{���M�1�e�f��N _r��º����QX**��裆��aPZ:4�H�~l���Z|Wp�h}�8���
����Fd�!���6[j� 6���!,�T���1Eu,
�e`���V�Ͱ&�0�q@BS�j�ߔ�W�Ct��\M�����E
4�ì�gCiY��ȡ2����F�\���xd���#�5��|\>�H��G=��� �t���Z>6%�K�jq �3��\::z�"Y�1�7FJ�Q����> ��zq�dV=�L]�*̴>��C/N�2C.?����Ͼ1s�z��3O6��Vk)O��M���dɅ"�Y���64:Qo�}Q�Ng_�G�24#����*r
�?�\ƝvQO�Ν,�-��lY}<�����L4v 9�'S�d�#F�<�ϊJܷ���0��!/���Ҽ�%���X�d+,���bܙ���������B>��}.O�+ѿ!嶄�� 5TEW�:�I��w�6AuvQI8��v�7���]�-�ِ���W����Z"�����*���t[L�}�Rlx��术�5G%ÿ-���)@��e+T������BQ)N����� d��(d�9#|�칧�]y��c�j�	��d������D�q����ķqD��o^tG!����c�s�?���&�E��HuX}��b�9/�(�)D�;7�=b��5�K�3e�ʨ:y�?��U��K�;<�=�}v���I�]�V���,��W��GU���^Ne�G��ǙD|�P9Ěn��]�i��}6��k�
�)���)�<��������!c���qOu�-:��n���R��Vn����s�'�ZRb�qul�l��P-�YQW�(�m_��5@���L�H"7�����$�'�F�q�� I삁��tP+�р���d4M3�u�����E�/��ju���hE���P)�U*\��X�j��WT�I�c��'̜��÷/�5'��}���w�jGEq�����N$ܵ��nh��t���/�-n�dL`B�Y�OS�r�]��k&�g�?������L�lMU/o5�!��8`��ɧ7CÜ`�|+��D>0��{��3޿@���1�q�����S�V1"ʥ�fC�L%�]Ů���5{�(g�yAw�9��D����dq�r�]�!#�3��`�M�Ԡ�j)��:K��xj!wü�SOT�z�ǂ/f3�2-��58-i���jM�Q�+�+�n�t|��a��Њj�Xg��H(��OQ���<�rţ[��X��)}a�&�M*l/0�����R0�=�c�d"[�=ȵm��&�3��⛲�I��¼���XZ���΂!�0s@4R�r�'� ��˯��!���ظB�v7�3����{3�d+��6q ������CŶ�Qh ��u�Tԁ��S���� t�3��q�2�h`t����K��\ц��])����y��K�F+燄��u�0�V��mv���z�WZ:M6wx<���Hn����;�G�
K�����. Uւ��&�|��WW茞�!ZE�4��]g�a�����і�D��7E�]7�τօ	o1j(���E��k�8�`[g�Z.�J�Ɩ�p�,K|߿d8��(�x��'/��M�)$Y�v%�Ȫg��I˛{�B|��L_�h�-�r&S�
k7����&5�b�wŹ4�����7�C�5�.���	mS�<u&�*D&�v�Hox��#�ܴ߹�x@�~�SHj�Z��޾�/��L��%��2��k2B�>�񸇂SC.ܐ��I��Q�g�
��@ev8Q8r�Q-H�6�����(d�"�u0:�q�0C�6��� "CR��_���@5�n�;��g|kZ�WX��$n�v~X�芹/nU����������"�3�j�`�n�㍌m��U#��|���x�:�3�E�����ŸI�����_���괈�5����E[��(x�k*�*�YY�x�N�`��)259ddi�=�b�7W	�/�F����L�R��0*-�m�1�4X87	���J��B�#b�X�Q.�`��;k�+�F��lbK�Q�NM+��3�����\]�-A�	jMӇ��a�8h�*A�!�C�L����0��{�e���|�J����pῃ��]� �n6���$T�;�k�N�,����f��0�P�ǝ��gޮ)������������'В�6))�:�}��[���X����2!0��3kKz�>�#�{\�dF�� ��UӼ���<B�'?���y|�M&;���;��F5ҁ�SZ��N
�&�k?�f���dD�ф&?�P��@("1[��X�� "s=���������j���bzd�\��2��%�~��?.	�]r.:� 9�S;��������+GB��A��b%a�ת��X�l3�n2��Y(���|���;�z�jI���X\���bM�S��j��"��s;{Te{�G�2�	���b��wO���Ů�ς@���1?�ew���q�q2S_���vԬ@q/z:̆��1����C��~�������������=}�Awj7���)��`-�F4��O�`��}�?r-��ؚ;-b������H��EBPDU����(�Y�tm{JO5)�e���s��t�ʨZ�-�.Q�Q�����v�Q>��Xtg�����) ��KY�����L�f��	9����p�p��I�-�/�3�@|`;�&�����Rw��U<�
\�h�/"
v�*�'y�q�����(��D�M��<QBJ�c���$���5��1p����@V�nOKe9�E4iB��p��^x1/Ŧ���UKY�.�g�b����e�a�]��
��H?K��D���0(g{�T�.�Xݣb$�vM�­}���F셩�3�������e<�͔s.^�cf1�����b�˾��k��O1t}�OKac��Kd�輲q�Csf�Q����}Ps�E��\r|u��
=[$��,v���f "h9(��l�7H	� �i�H�9Do��M��^.A��t))oq��{�"�ix6v~eNCT(H�V�������r����J�e�5��h�`:{ga4+_�h��o��,Ž_�v�������>{������"�h���Y���@�s�v�Y�W���d_]9������.��~���"$q�eٓ�Q�ݯs�gU���d�-�y��O�CYF��)�9�3.��:��"٥��Ԇ�t�w�E�Ikj��k�w'� �� "����M��#�b��ĭ`X�=~nQ3/��H>�Z�!-��@�Y�_�����|�lO�*��6f�N�",pV	��L��C��3�Vg��qy����S�Nb�j
k��y�v������za<�VM�0�X���<!(7�'��Vg�\Rkܶw�{�,�sH�*��	��\D7.K` ��1�c� `.��p*/N��',�b$�^����#�v�=EMb,�$��͔C��a�����NfH�S�L�2SJ�@����A����]s���"�P��k�V����H}�0{7�~����q~a��MQv�ؠn���p��|^U�iJ�m</p�݃�:�S�ZG㯚�2��Ȏ��xtJ��r�k��|zJ�8�;9���}º��YVX�B����w@f��0d�^?��rS�V�yÌ���X�e��_����oZn�H�=n,�͸�.Z ];��j-�{8�����c����:`Y��Ǣ|NG	��Dq��?��}}%���;�����uׂ�eNA�������a�Q���η�f���Iڀ����;�Vo (�u����5��J�R$��/⳸B�6�3N�Q�Kz�ac��k.ؾ����0R�FG���k�� �C��}�y*W���uJ�2lL��{3I[�^(g�N�K�I�hŏ�O	uUC}��*j�9b:E��]�>����pAX軁o�ي���(ȹ��s6`��/�EI�/��)_<���yOcA�'<|�k8�3�<�:۰ANVNQ���͟uL7pܥK`���@.��_Yi\`�N*	S����@�����M�����!�c�	!3~��J���枠��V���:��D`�
�ʮ���=O�ޝ�+p�x5C����{���Q��.���c��{��t�J��Wk!ɣ�����b.4�$�+6��S����B\�[�vC�r�MmS�lu�6�^&̼����-p2��Q�����D�F�����u�͕ߍD��]�HX�o���z�A����gB���[�*��1�O�v�H�����%����t����w���C���@x-��=�p���#�AA���c�./ �^��o4ԙ��YQL�6�>c-��̻v7>�΢fU���g�M5T���r�c�b��g��0t��b�K.�!P�!���[hx�=�⺤��v��#:O�ZK�&����ǘ�������n�!]G�4,�I8��Nߌ?_�]���)Pg�lv*�X;(�����[�i���঵�E��hr�tr^�=���a��S������Y�[��'_�\Ą�&��F�R`�gY'�����\�Ͳ��y��!��b�T����ɉ�������2?�,P�(A��+��by@	��=��	�ݭ��,��q�Qq(B�������x�1h;��#�2X4>�����2�����i�ܩ��q�:v4�]
�%q�G�� )A9�w���Uc��T����_��Fhz	�*S�y��qh�H�)���<-�-��)&9��z��p�?JNV,��55�r'!P��.�|�m(N-�q+hK�z^�I�^(�� �D�%���{�[
a���n
B�6\���u���Sg\��)3��샀�h�{��&v\�`/\x,�N�7�}����GCvG�!?Yq&��%�@���Iߘ�`y�oOp�G)�ƃ�,v��$R}PJ�K��9�i�>Ȃ_Zq����=`_�}r���O�</�ە~��47�}�t��8<&8~�SׇmWe�L.�;3c�c�g-F)�AcT/�d[8��3)p�K�'�+���EQ�Ji�.H�*�%\�B#P;�a�����DI�HP��hЪՓ�K�ۦ0q�El+�`�p���D�p����8%�[�gK��ig7�����Q��ں�[�j���;QWψ�YB&��=�e桸��U~��.O�c�����8��]�;i�p_F�[�I����b�j́;�` %��'��t��W�Ǟ�좼bL��g�s��2$�!��\��,��9�6����}_�I>tD�h�ROr�\u����+��� R��b�r���m����-}c ���e���-�=��#�r�!����JMZ�)Ϳ�S��T���A_���$�}��2QUy�
;�
W�����m����������$Y��,�c���e����F\8�Uk'i�?��Y�\|a��	�0qK����K�Jc-��l�����$B�D�E�a�Z.�X�Ru�A�b��Xw|A-ɍ��%�$rRs��%1JX�ˇ�������;�P�ߑX��b0ЃV��땉���T�p��Qo�y6w��$� A=(����Hwն�U��k���%�GT��U9x������4[DK��8(	����S���J�g+Ԣ�=ئ��B�[i-ar�O�#�=�~W�wY�?ˋ9��s����`W?Q��s:��j{���ȗ|�w��4���ܕ�|����|���T����)vPpR�6�r��K1O�,�{�������S#[W�m|����0��O�K���2��}9�,0���n�Y�������7р��E΍��8�}�����E�s_�wd�<�;e{|��0�A����W�jY��G�4�p%�{��ne�.��CmP��*�h=�8���f�p���i�`��8A���f$ɷ�M�d�o�2Ȅ�A���}moMm5�~���7-Ws��Z\e���:(�20�e��"��U�����x��r?�}�A���SJ�!�;����d�\a`��]7/��5�t�~ }��k������l�	C	 Z 0�5AICcM�������ei| �I��B"#�`�A���qp=��ĉ�!��qܙ~9\�]G v"�����+�SÙ`{��=�c�_�X�����ץ�����Ɔ�6�Y5�uV�T�<��va���j��`A�]�{��G)e6|9C*��x#�����k�|���%ָ���/���>W_P<�-�h�5<9�/����:�4�?k�r���cgf�u5e^�?ŷ��  t���h����]�i�m��&o��q���Z�+V����5������W�XD�4��*�>^r�ζ'#t��D}VYa;>�'���^�@�#�#͗2���͝��j���F�X��h+X�&ζј���@�Pߒ�,�s;G�So��GG%+]�fV���6�R�:�/޽��X�� ���J먺��j�b-����5-�z�t�(�<6��8�^��	*<!�Xx�L��E�s��