��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�KW�UHսm0{�K����ّ�����pz_o AHs�=��r���]���J� �o���1�(�����D�[����*��*m
;�{�H�i�H
����W���� v��Fo�:]Vb�"WB>�`�*0�=|d���-e�X���������liz�ٶ�1V����U�$0Xm����OV_!���&܉�R��.K�ӥ�U��S�a�;{:ŕx=b��1i,��N�Jp
yg��N�/�:�x��E=|}`{V��o~w��c��V�9��c�IK����r}�F�ظ&�QM���fș�,斐�k3iQ���n��?���q�X�A���o���9����5�i9WtJvd�J m6�@�
�9	8$����&\���,��S���^�_ѭd��W�+�{��c�~-��*�#���,r�;�(�돋�'��v/!*�����i2%ĪkN�$��3Vgva`v�p���H�z�y�J'�ȉ��+o����)!G�*��FΫ�
��Iz�����W�?!���������zU2��4�H�K�Ѕ�?�	j|�{�У����uZ��VsXD��]�6y��?A���tٚ�1W�6��?��>� Q�C�0�E������r
!>�O��D��6�Y�~/.�1�t*��O\J���T1�a�&���n����;&�q�r��_�6��G��K Я��������z2���T��J�V�>\�P��t�Sc�vh�����e�Z
�7��Л�S}���+:�X���{���7��u;�Ϻ7Ȉ��#b��M6{���V{�oE���FH�o�2�ĿP���v�`� u��I��ܮ6�4��4���[KݷEl���G�sn�`Ф����)�W�4��J�-�� Š��ᯠ/���P0�O�ޥ�d��v_>k.vBz��*q �3و�z�R{���Ļ�~�FȎ�IH���wb$V�u�-��C�z5�}�&�<I�c���騅��U�PP��Fq��u(^'ǹr��Nyj8���I��r���O�i�����c�r�~n��p]�z1�1p��;�O1�.y.uΣ(����r�ܽ�%�1�3/�z\�5=6v��y���� �dw1x���ȧr�!��h��[߬x= SR�8��� )H��.�d�-�V��/�u�X���|�@{aG��$��ؤ8��t΃3֙(YF,�gv�K^$\�q�9@���5�<��p�bg7MŞɼj� �#ɑ�8�S�<q�R=�;�{^M] ��~mycK��+��r�
z1�W�g�� �X�1��>{�}J�Bvy?��A����\�� %��X[R6b+�s���E����Et:z�7�]�B	#�D�x�EO�NզOƣ@��MB�Pc�呁���^����T1���wF=��
E@�ᨃc]ne��Db�z};	��}��T�?��'�-H���A�<8�S�\C��E��b�R���<�� ��$	L�l;����<?К��[eԥRhz�9Q\Րd|lO�Gs��+�����}�D�Ea̼��mb�q��3}T�g�k "��,��g��<э�|���4���s�5��p�X�	���fL,Qf����&�b���콁�<�O��H��|���m��ԭ�<b�~����;��ߙ��k�.�?��{��k���� e%X�g<�7u�٩�ԁ�O�l����Ǌ���) c2�Z��զ�Z1����톺/�PU�E+�榚7�<�]�@�`̺��[s�Ҽ.H��^ꌬ�VH�����
�u�|�d����u�����J��o�f'?Uߴ�c2 �mO&���땧\�Gy�[����:������ޱ�0Yt�dv��&�RҺ�����X��&Ŀb��(v�S�#�9D7^�r�U
�GGTE57X�9}�-g�@��=�(A�ʹ�g�D.S=�	٢�/@EG���{uh5*G�&f h\"!#ـa�]ye�]|Wج����� �<}Z�W�>����g���mb'�@
�U�Δ�r'���_�2�I�Ȣ����X`�;T�,{�O��Sl�s��r^�|�]���"�lb�{��/�ǯ#��~�>�ۘ�0�F�3�1�����6(�Dҍ�Sl�l��t�Uz�X��q�M��Ul ���X��	��8�`�e���n���F�oao��"�l�~�s��9�X����I>vQqL)�_�(���Bp����v�&��s�Uݐ`��B�k������k���
���Hb�}��, Ɓ���¦���V��,ދ�4�2��G�}&�C���WRU����8gA��3�M�R����^�S�(��#6���㪱V�ͨN=x][=��%B�i�����:�֫��V�g~ơf�����v�춌��|  �y�J'�svc@V�6Y�M5�e�|��{/4L$^I�5AH�9f�q-eJ�u 1�тv"P"Bݧ�LvO�{����h�����F����1���5���G^��/vU im��4s�eD>�K���-Ӓ2idå��j��KQ<I�t�:�؉;;���5��8+��'�"=�O��ԩI��0ɻ�Wm�[���"���[
K}��E�+�7�Vk`�����h!ŏ>�m!��l�ɟʋ��h��k������������E^��-S]�X�K�����*��:M���c�J���3��h�;2�Q`O=�c��qa�ޣ.�Nbe��"ݦ�N�S3z��]�Q ����9a3�+W�F׊+�z��`2���&��1߬��o2_��X�	����_�!������'�r�X?2��)��f�`V��0HB��ɱ�G�,���ʊ��q���+hh�N�����j� �O��e/����?Mk��+'�����3�PM�I)'=4}����i��[�K�\g�Iz����>������$�ϭ0)��9qa�����C;+�1N���N@rh0�!.6lZ�I�
�1�����%<���{��rc���u��R��r!�o�K?�q��i�U������j��=�BNp3c�iFaQ��,�IiX��Av�@A')Io�p�1����������*TA3������V���YqwP!����`��'�͜�����{b�wp���1�,�8z\�B��N��	�o�".?�|�=`�z�C��thS�k���.�Θ��MW�p����V����j�����/�ŤC�F\��a˪:�V�*��$\�+��o5�/V���t��.��q��g�A��b�b��B;(P�:� oT�~4B8h�;8��Q��v"@	�a�
�q���g� P3�?������F?�N�*����v�f�9�� �#n��v���Q�p�	a3o�b\��~4��7�ua��.^C6#E�٠F�E���K�0�/��CiB��VY9����U���)�v��M<:c�ьi��+�������7}|o��C�\��|0>ʍ�~�<��������~�E�X�xp�e�+x��tjr*n]=���r�9�nM�h�*`�ڑ���\�+��u:o��q�e:�b�����5��4��=V;�&�=�I2����]h�Af5�����ק�*����{��^s��@�=�sf)���#�c�r�r���I����(�1��`%Y��ŉ*�?�Y�<�N�cOe�y�^O}�bk�̂�LI�Mh$1~�Q$��%V㥵ye0o��ۯe�p��L��'?�Wy�gX<�K"�uD�B=l��Rv�^H�I�� O�~=9 ��w��uL�����</{��1q%i���<�$L��Y�R�t�f�I2��_(a�.��-LŪlf��9����Y���ǟ ��m�1�Ɩ�B���x3���(̮����� ����7��:y1�p��ȴe��+nu�z����݆��fN�y��%�,i׺��������Y�'���6��4ڄm,:��Rz{��tܒ���Ȋ9����4����pq���4D�|���u̪�'�E�'؊e�c{Uvp��wI|j�Ӷ ���vZ�j�9��K��Z���͹9���~Q��?pؗ����R��D���[�]|�����
��2�4}E��oﮎ� ���E5r��,�L4�-��IN���
��	P���>׳m�a�-N1;Pf#,C;��s�g�E	�W���W�@/�i�(�dX
�m3�$��k7�&��A��v�Ea�[8W���̆@K47Gŧ@U��"� >T�Z��E��� ��+kgmz���� �ȲG��� ����Ғ��ѕ`g��.�E�#��=����m���1վ:���<�@���
�ޠ[%D��A��b�ȱ�,���?�҅�J.�����Ԓ�Wq��%1���7*� �8d�Y��-��dh���5GS[��G���F�r*�p�C��GjN��U�������S�{�9M��(�u�����J.!.w��I㢅�Z�3F�M����̤��T@�6G���}h��*�M���Vyd~N�*CKΚ�>�a$���Ř(@��i{��㽥�_��������;q/��Z�U>�ӎ��Y+-8 G1NGZ��I��S՘]ljR~똈(�5܈�3{��8q�t��{A�K���sC��~Q��D"`,�ě_|�C�x������(�ް�H�Eك��8�8G�7}F�ONn½����������� 2�C���WN7�
{c6���Қ>�*̦��x�4�j������P�J��3�v�]���	0�[�%�tG�G��s��[��|'������i�S�4!���D�\i��;�x̗�ۣ�	h�{I����������)�Kg�T�����"���yUk�]��{���x�������ʵ����TQ0:l�b�j�t��Y4)x힞�1��Cz��裠�AN�� }�$d�Դ6��_SA�>��_�����s	��^�,4���'o�����!�P6��~9Z�����"��	E���:2`��M���HQp�|�~�8��.�>&>2�u�Q�7*_ɗ7��aM�,�{q���z��?[�q¯}��0&�6Z��a2B�7����;���>����!��F,��7�� �z3i�g*cX	�n�P��%/�i��`�����T�ip��<&�#&�S��6��;�<��L$'���I��:jma�DV�ݻ�xW�g���Q��ǚ}�H7�B/S6��㖓��p���F�3dl����r����I�lU�,2�y_`�#���T�Į�{N����59�2TPÿN�A�7��	��בo�7�)Mv�*/JֿBD�:2�����w�P*Dڗi$���l�#���s�8HN���z�ӮOQn�������y��jE���c���B�oO�LT {�U������[?y]�����&p�`*m+O�pf)`��C�YkM3]�J�ޖN�V=�����ʎ��>�A��,��Y��DQ�*9?o�Gd���J�1|���k���FM�i��~[�En��Ib�@���>���%gl�A�A$Rz͛8�?�E{�pU@r�j�|J�,y#��ǌ�[�5vG�v��Y�5Č�odv��ň��ؓ�@*EW��q� ��h�`P؀��T׺���n�*�=0t��;�B��hO���H�L4��Nt�"��eU�{iq�R���H�9�e����t�n��*�~E��(^�^�z��&��33ޣd����~.Eޘ��)[oAf���t U�"����f3.1�=�f39��V���l�)NX��"{K��a���	��/�8�6����<v���aHH-+Z���y�7��+5�9��۠�)?�[��V��ڶ�/إ;��X'Y"Ub���8���Gz���ܡZ��U2�L�*�e��P�a�$6��j�J8Q�،.���~>rX�9�I���Y��Ai8_�AF�O %��b�����9t��k��x*ɠ�4���X���e����;RG`M�2��f
k|�p=ŷjcr#�{C�_Zf��s��5��, |!��o�7;rG�aY�T���M�Q2�E��X/l��?��Ziy����+[]:?A�LG�_a̿t<��=��%/i�@2���b$=��
���!��4Е����l������g%���rw��I�l�B`��I�x\��HłZ~�J�}���B���
 ���@��}U�G�w�f�
Z�~����v����[<$`r���^y����͍�O�@/�i��(8�d]��h�޼@d���^�7�/!��E��S�y(����n�[�\t~@�fB�a 7 �)��t2��h���C�swAs.m�9K;ϸ�'��L�}i��Y��Q-��w�0�H���:�� t�`�~���ȥ��~P�ԇ/�O�ӊ��ȯsa-ُ���q�6����,2��]`vu���$=���%����0�DH�?�b�Gs��5����y�DC���i���(M�}��-BPu
5��b���Q�-�8	�G��F���kSЋ��{��G�	
�M�/�K�Y�Ѭ�~��uq�˚S�]����&�.�^l�m��o�0y� YxŶ����^����6z�掺��15����2�V�ďl�3.W���ҧ�:�/	�p���V�A�����o���:y�H�o���J�s7`�焱y�T���	��� 9^���0uj_�������N��8/p�
��{q=槂�P%{��[MXfqg�,��d��̡�t��r��u�� [>�¼� �-�8��yu�LI6�EjT���h8�Q�m����� �	x�!:Z��,Ec<Y��ݣ&e���u�`�������0+�Z��Ӿ�IӖ�"+����\���xH�)$fX�����������i���'f��C��s�(�Ot�� `��g�1�+B� |�b�u)D�y7��EH�)���ֈ�{�~���s>��S?�5O���N@�v��Ϝ�G�͢5r;�����2f����:�GA����r_+m^�$@)�ׂ�MF�<�h*�+!�eZ�z�Y@�f��A�6�	���"�	=[�>[֟݌?�oy�?��Jy�"��I��N��z
bnD?���@x��Dߩ򺳁?I�k��M��e���F{��ۂhb5���g}��%�:q�O��?%\E�y�����P��yB)`�Ъ�h4�5 ���,*�j�A��J��V�ǳ�L��~��)T�o.`�-?؃���F۝��y�$��iS�]��K���ʗ� �Y;QPm�z4���f�F0���2��f���c)Kzb�XY�J�~�$����H��?�n���f�嘺Ir��s�����ޡlUp)�n��ډ�%�"�IɒSp�K�x�����5�Ӧ���XIxWx2`lc��ΞQV1�Ca3�긳:��p��9���� OMf�����1�!Nc�J���)���Źwy<\�ڱ7�� ;�Nݼ���,�n����!g����􈕢����݁<�j!ӋaɈ�c-��~��(B;@ɷ�Z����u�郑f_R��������gL#��wl��~�����@��W@�8��70T���~�_ U�������Mwf������H���O���;����Q�c�p���*"oq�4�6���Е�B�E��aEW�Ǹ"����h�ﰶ�y%��# a���0������G+=�Be7��y�z��d���$�f6@c�︓��9ML��L��ڀW����^�K�iŷ�6��Yc�X����HLE�Ek�0c�f6*��j���WH��]�<��گ�3^9�Q�;��[GQ*��헞X�)�6�r�8)���v��PeY�s)�މ����������\j����e�r�eU'�9�X4���QY\@&S��Y{y�8v�K�^"$f<�ɠ��̷8�U��)�aT  ���eE-��^��:�����sO=(��G���	��10|������!����R��_5t�)��nz����٭1J�r�Iu�
��Y�r�E��+�A�(���5}��m���pQ^�A�B��z0���U��R�vzoơ�v#�2�Tw�#����	��~��&��c���d����(�l��VLk^Јk�ίY��)B���[l���������R��U�=��%��n�5��ŠD"��l�9A�	�|���s�d�2N�
�B�;'2�+h,����Añ���`��D"'IT]���0X$F���)3#3�@�*5'�T���3�
�y�O�YM{�=��8�rO?u�/�:t���顯��WP1�U�F2���l�����fX�Ռ �&�Į��0t���{
�K0���-a��3,SF�u�E܁�4���)�%s����(�����H����+N675�4ٙ�d'�t;�LĚI�o�;+)8r��t3w)bM�����.&CLxѣ��wz`��(�"�9�{�
��@-7�n��O0���5�!�ߠֵ3�}<�0�H�P?b�����@S�>g���k�2��~׹zi��ț���U�}���m�9�$�����j¥$�]��]��~�{��&B���)�hmܠaIw�9�"t��3���Z���Z�^l�^���;��}5���#��Q��u6�dl���A�P"w�	)V���r����0o
�&�%�~�
��L��ڼ7�$�j^����a��6�4l����&�{wRW���jM����M�Fҥ������`�H�ج4�h?����2��%���)�G2H�zѾhJu��Q�:�7�]{v@�6}zc* �� ��>�� ?K��N���q��R�`\)�1�6,Oݬ�!�U�J�Xrgr�D�/������j�o�;���"B���x��{���.1�k?:&����2�=KV���v�E٫#w��];���xw��E��PQ���7�a�(��J����~�(Mg���}�Ւ�@�>�2�Cm�uTp,��O�kGL4�6HZ:���O*��]���.��).�2����A|�K�:�_MH��뭢������^���1�;^�0%�T0�F9$���lp���I�#ތ���
;=( ��H{.!�ȼ�0�S9��/5��f���T;h����������UkʭUf7�%o>��l��{%�C���Q��}�w,ףVW�R )d�����K?�Vt�k+=��zf�|;N+j^���VW���rϢ���s�S%���9<�|�2�>�����PB��$�I��]2����ϧ�X����O`θt!j��J�
�/�IB�܏�.������3,�������A�+��x�=���~]%�I[T��複��{_�kݷa�����@](Y�O,ז��$��^w/��@J���J����b߻�6HZ�tF�B�$}�q�w�����<��9�����4�J����Z^V�tgT9f��Z�ݸ���&�!g_�J����鱚ѪAל�هY�G
KY����p��� �G��W�b�%���t�8j�����ص=THaل [\8���LCŲ��g*�>�j��P��%��1JW੆FZ�����Uz����Bz�?56��
()���׊���h�$LϦB�mq�G#YD���e�S���P����vq�s���Q
~psٚ?�f��_E{�_�?�G�=�C�Ԉ�������c��f<.��="v~/��|�N��p��͘��M��jy���ie��-S[��������nz��4a�X�~���=�d%�����N�XB8���A�ē�E;xa��X�:���6�{�sjƍ���(¿���m����d�O}4�wÏ��]xƥ���&��eZ6���'w�3�q���~٭���3cs�y����!oe��\�Y���We�Zb�a�,�*U���ؠ*�>�N��a�K������� v�@���g������XWO[�w���D2�$��0��__'����l����z�=	���'�	���a���b���t�3�|���7��m46OV�!��5C��bC�3�n�\�;�yf%%w���F����Bui�m����Ӵ�EO��7����U4�5� 2�kTs�>:_3��B0C��T�ФV��%�΋��]T|/�5�����a�r$	�D7b�,��r���E�6 �B�u�y�@)Kјb42t@ڮh���<Q�P�z����a��t�!��Ons�DޮQK���;�g�^`1Pò�ok,D����د	>�=��1��\��\ٲd�e��������G3�K�C��5�(�*���L:�|�-?���1�{3G��8�9�V���1ɵ�chO%y�b�U8(��oU�^�Y�[xݓ���|��K�;���S�jm���--�k�d�k1�x�D;�W�*�A�ea�ʤ�A�Z�	6����*) �9�G�9n���Wº���h郙�0���Zi7mv|���n�X�nf\�:10{Y~��ы(W<�����/ �6�ء'w�!X�Ιi6��B��{6�;�.�}�`��Q{��y��."�kmT7�aWp��H%@��q�E3���������$r�؅,1����\�pt��(f�F:>�p��|D��`ɚh��N{��	�5NRTTA���D���g5Lًv�v4���������N�%�O]o��'i���y^t�L�������(2a��fd&0���\l�,�H��3i��-��$����M�_ݍZ]�@��T��}��J4![h�	[0&cؤձ�qq����d���:"���;. ����D3 �2`H��Cs8�����zm�9墌�L~;�2ȁ#�vT���07Y�Jø~�T��Z����]�Tg�Հ �ґ�k	�nGi�����k��p|7Z��n�}�OnYٰ�v:�w)*s��Y��t����`F�
�����hK���('߄Ε�K�tf���B:D��,?~̪�*�F�X-ڏ;3���*?�=���\�n�t*��1��[����)���{l�*ح=/��7��W��V"'"�`35F�6X,|�*�e���/6�<�h�w�tWi!?cA��$��B����4��h;��e-��֞�����M��hr�#ɐl�l��w}�Nm՟�'h?�];>W��|����ћ�e�<�v�q��Q��p��(��!�Ȫc�ϡ�.VD?OĤ�sU^�����ך��b��.d �P����U~�����d;� �db�!����h��E�p�.�A���'�L%�Ò���x��Y�~�J?�.`��^l}���4㊈�1&��
�p�_D��f��Yi�ZJS7]F��]IN�&�oZ�RŦu�X��d�Z͜�w�5�;�~�5����8~�:�$�:!�]"Ok;D
o=(� MT�	О���l��z��OM�:<�Ѝ�nÞ����gH*g���932 _]G.2�儆�Y�0ʫ��(r�z屮;)�+�x=*=:��6��Ie�����<���^S����۰^��8�՗G.�@�)�lza�|_᧥���e��A�t�|ȍ1�V�>�7뢦"jO��MCm[�ݥF���k�	G|	jh(W��j/�ީ�1�馶zY���������Z�MD!�����c��ʿd�)�jN�1�mjYU�]ȥg�i#"u�3�V�!dK�	y��M��<����9C0�F�?��Ν��	%�$����3�G0�c����+ُ>��L�L|� v	yr�1�s��w�j����`B6��.6׭�+�v��[�g���ci�����¹*����+��l��»��ְ9�oR�?�k����L�j� ��	
	��d�K��(�CƤߑ�!��Kx�I�����`P��\�>�e%��!$��}�I5A���X�/�X`-jU�e���F����{�	��\�$1s�����S�.hV0���[��b��r'�2B����K�nw0�U9���F�S�I��4j�Y�~�Ӓ}��P=��
���{U@�B(O���3�z@��n��D�T�XkI��s�QC��;so]sDX�D�j���0�o��
W{`w�F��p���}^y��>>a�Uu��_ȵ
��@�\@�����L��Б��[ё�-��ߎ�ƞ�0P���N�\XJ��7�g��?��+�W/���g���7��}4s�fA=�9^�7
'��<��*��#���x��~0�kH�;���a��/U�q��5m{|u�;+��_:�x4Ny�EH�;+eh��ކm/�����}�a�W�4�	m\�&��6�w�>�����!�`��l��$Vp1>�
�_G�Q�$_4�h��Q��KS/��V��z���ӣ��#2q��m�Ā����[�ʟ� �Ya��;�$��1|�Aqt�b#tٰ�)+u�.k�d�c�%�-��c<'�4�����D�{#{�-��	�0F�~.�B��b�6��x#r�H�<��Y�D	T�<.F��6d7n�6�����j`����K�H ?�ZY>�c��\f�)Ϫ�xJ�{�s@�U�@z�#�����#� S*�7�gn�"�w�q�����T���������M�od
����C�-����N�:�ȧ�p-���l��ŋ&�2�Z�[�E��tP"W��j�&܋�U��Mf
�����&I7˫��j1��D�1�w_��O�q��Sc6��ف8�/X_��eQՈ��ő���p8�0����D��j�{۽w�yċ�����"K1��P��Z]��C@���G�G�ƠiR��z>��R�Ge�����q *ϕ�����Qa��� �Ot��D
"0K<7�Ggq���:�'A��-(q�ۏu����r��l:��c�E�Ր$"��:2�jw��5Z;�Y�e�:�]0���q���Dq��i���o��G���|�p�A�0ȩ�2��
;-<�4�-;_{�: �fc�r�噜2.�GA&߆��7�'���B����kBC)��ꡑ�-gw)�@ ^̀��HN���o����:�4����e�3O�F�(E�����6v2v���j�7�9 ���o�ɰ�6;/�`��@�GQ �q��u�m���r�1�^_�h�E��%S�஫޶�#�S$�o�n�|NM�������x	]S�&����5�?��/ȸ���!�_n�u~�,�q].��F\��oB�D���9��9��(\xCu�����d��Pr2Y���L|8������/�M٤S�I�?���{ s���/2�?Upڳ@��CRrw���L�=R��K'��fN3�|�&����o	�]��T��6���H��b��ƦjCԵ$*���G� ��D0��/S(vxщ���c�����R�3ȁ�q�a�l��^P��m���"���2���J
ߝ�+���aoYә�ī�$g�g���Q�����x��ȶT�\�v��s�3��X�	��$H?IP� T��?��d�:�ƣk3���J��4�S���ǉ�Q�����|��/�%�٣+�?��q�6�ك�`�*X�� g��c�׺:'�H�]�N�>�*�U���[��y-굃τ�HV�V��U?�Q0*S��t	���K�Vd��y&we��'��H�p�Q`V3W3�{D�:�͗�G��������ACqH�^0x���BY_@8`z�K�j���&�ҁh�ZvN���%6e�x��s����>���^u[�܁p�����BEa��:�+sN-�a�������n��V���A�]O����'b�'�� �B�VSM��)<ɜK��26���/H���ֻ`��;@��Ŭ��||kAw��\��������L�2�Z\���bTt;��)����q�F	b>mr3����%X�����[�H����GQ�j�&Fr��G�ճ�k8��~�:9q�X-�6�A;u�b[%7pEsS�=;�-Y����t�����\�a�`(Pľ���L����Wrp��4<.b��1ߺ�׀a����q��3�2�}���bo�ٖ�����2g�<�<��.-��=���M�5^k,�.��wq�9����T���J���5��(-WSXg��L��[����K)y�Qe�=C)��̆d������ �{+���J�8&���`�ՙ��'nB��b��(��=�}t�j���iyM���O]�u�[p�y"%6U<ᶧ'��H��ō��({t�ژr�(�~�@2��ށ�r�`��O�I��lQ+g񛖕�k����d��ar���K�?}�@�5�b��&�>��L�kW���bWdB�3�\-"�{.�{{[ӥy��Y��zf(�0�a��6���0��Q.�a~���|���s$%LI�Ns����%�4%NN��>Tz~�Y�w["dPLO��7D@�a|�w'L����c�����K�7�DD\��0N{���xUoi��
���ve5t��f��^"<QXA0�ũ�k�^*����˻�7i�	�C�lDғ�M�7!��2�o�|���Sa���.�%�����,玒Aj�'�.N�������I<F�������[�H���?$A�R�����Gfb����}��j�f���a��֠t �W��UͲ��%r7�*L'=8<He�6���>h�]��&�����T��	 �h΄��~ �p.�_�tMj��Xx$�����^Rb�~-A�6ϖ�����V6��3cנ(���H��锲W5;��R����!���>���i�'h��?&�!{� �&�����p[E��ٞ��ADN�����5�E�0ka��>2L�����������3�g�Z�G,W���˵e5.FjDە�^��ٰZ����BrX�Ϳp�s�+q� AOg7���"G�K�l2,�y��%'��o�1]�jt��ط�e�K��2���� �Q2$GR�O�\G���A��:����Ǚ���ǳ���'��N���a�x�y*.*��G�dI�EM���B�ˊ&O�>Cm�R`�n�t3�I���S;��|̴*&�H��� �a��\9�֧�扔L�g�?٢	Zސ�D�S3ڶ>6�Ÿֺ�C�A�5~�ߦB�X�����Ƭ����C�Z!rN�P��@AT��j�:�|��+_t\蝓��aN�2��ɒ�q��-z�� �R�k\����E��zq:��g&>�O,��Z�ʚ�로��W-z��,��k���6���F� GwxN�sY��2���*���C�������V�� ��i 2\���v�OA@��Ş�K�XɄ1���h1g����@��7��K#�(+:8�c;��-�����\�S,(b�jK���a���v���|�{�2��Y.��o�ɖ��U�2>v�OG���/H��G�H/p�w*A��f���*�A���@�����-1?���p����&Q$�S+qٽ�(��|!������.�&�N�,�Js���inT�_2�јN����5h=;�2D��{�+m��+E��֎=��i�߂^���v���e�j��|o��(��8�Z�J%�g\EUaD�hP����n���|^u4̼�Hٞ>����=\���3�����ɷ9 ;�Iʌ�R���F*ӷ�2��.΂����iM}����%�/:�d|�9����imT���Z�Q��K��S��o
�Ҝz���)8��7c����5XÂ�&�h_�Z���8x��r��jɪb��/���k�a��a�T��`n���K�p'`���I�!��~���J(��A�<��Ib��䗴!Ao���X[2	ml�ig���&�dH�+���*[~x0O�E'X�