��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾���b������o��ǅ�}|XBi�v���Ĭ���DT�7ׁ��X/����J�(2h�sݤ��E��]u/��Jb;�A�����G��}�n�:9YQlX�,��K��:i��d�����I[��1���DQ�!���p6Щ�§���Mr�<`����=��Ece������"����"���]��h��ɱ3�� ��T��S%.q�_��u�-�F� L� �E�t��)��0��{{����cpA��k��z|j�9�� c_�y��j��}4�F~��U�·H��x�pV��i�߃?Lu�v'W�_nb�.�a�SL�}�����&G>�c�
;������6`Cz�h�,Co��ΐ�7|'�o��ÖF�[;��'�?v��2��^ ������(�(��~ܣc���<b6[�X�?����a|]b���8�\�]&~��içrq�G?��w��e��X�6&�Mz�X�R�87��E�kw����
3W0U诵�6^���υ�����]p�G��HI�ip�{}�U����҂��Y�R�ѿ����lk TBM*����
�3��4UZ�}KA��!o�'��lCv]n��~� ��R�=�
T��z��x�D=�
�~�ozڙ�Y�<���a'�Ϩ�t��Ү`)}"%�w8�;7�<�}�R�wB)��٘@Θn�.y���L�%M�x��`s�7 :�c��/d~s�8���*}D�+�z�QeI[����&���5oz<���;8��
M>�UQ�ܙ'1����a3�:0O����Dw�n"��N24A��?`4)���������_t�TR)Y�`��h� q&"U�P7=��vq�N������S�&�������������<K�^�j�)ƃ*{c�TXN�\�;��T�p7���o�	�c��̸�n���R'_�|�|�7��ʹ�:p����R�U/���~v|!�պ,/cpa"�}p���ӻ�̱b%`&��/����c��vR���a��������V�,w�{�*1�U�i=��o��i�pҩ>��	��!bъ��hrE��ݼ�v���^��޺,�����0@ɔ�!��?�AAr��SU!~aˊ�nWG'�AC�M悄q��g�KV�UB���G,\q�ud�Im�Y��J�E�޴9�h�¶\��iKl��F�!o��~�X��SA�Dw-�:O�Ve� �.*8QdM�g�ɹ�ⷳCۃ	h64����C�e<U|����m�wkLt��a~��K����[�T�"k��/�=D�au����Ҿ�����I1��c�7�)�\�Y��/D �2Uh�_x�@O�g5Tþ 
�A�YZr���'����Qu�0I'��eU��F�e�E)+��o�F���Ķ�'��O����d"��Œ�,d�ιS}�ϐ�W��dۛ3����D����ñ6�#�ۏ~5%��ƍ�*�����|(����#>�ŝh$H#&Pk44@�w�s`����& pc��PitA26�7��6��1�����g(酀�����7Jg\��ˋZL�hb_���x9�/�4�eUbv9R�[��d!G�����S���0�VH2��O�@��Ӭ�	_���S9~�j��h!'W��&I�^�q6j�p5�
�ï#��v�
����Ԅp5G�>�l�o�,aJhK��se�WNTJ[�)���8����7S�����B� �5�K���q�S�V G%^�S�n�za'hc�,KK�vD����|�d}�
�%J)fQv`�oo:�Z�@da����9q2�|/�Qpe{uӤ�	��)��r�T���{�B��-����0�16�	�,��X�u�W����,�}U��AU(�Sv^F]l> G��7De�ٿM�I���'& ��	z���-EW�0UUn�oT��~6D�,/��O��S�#4�\�Z$�A,��2R�ZZ~��/϶�~��~G]#������i<�ϫض[��yfYC�V����LP��P���W�l��6������u��+��\�_��&yʂ�3cGO���P�(1X��q��+#=}��e#�9F���\_3*)�|A����%0E�gS�m���`��b�����C��`����C%�������� Z|�s�V9�6�8Σ�N���ݣS�僔��)y��`�>-,@Ն����18��L���}7 ���t>q�����|4����'�=��e�A�r6����KQ�Ю���F[��'��'�>���e�̓���������g�,*����ITe\�9t�f�n�����p1d�g<�(t<<�,�2�κ�w�!�ٙ�'l~�������)���i�dՐnc���o�J$��o��m���g��ҷ����/��܃�+J|g$�T!��@N!����; |%��ghDs0]ʻp$.O�=[�7a�ܼ��v?���-7ۢ�z6�vN|�s�ƣ�2yq�i|�~Se$��T.�ά�帩I�Ti�h� B:�c���`��_(��P-�zTH�C�q5��@�8mv��F��@_�A;���<�˞C�D�3�zB�F�6Q*���͋�Q�vt�ʲQɊŲڏ���$g���ݚ��b�/�tCn��D{�}�@�e[qCc�Ӕ?'�ɶ]�e���f����Zm j���-x��2X�]X���ʕ��vX�f$gyV1)���lI��Wũ=�s�-��~��F����t��:#�sU����7"z_��\�D��'1��TA�����q��z	 ؟��R�/�46;����,_E�zcTU��c��ݣ�\tkԱ�X�%<��~Xg�{/�^��+�g$�f\�q4^��h��e�^�|�@���q~p#
氤� ྼ�~f��!]�� �	���9,==�{��[�$�k��R�6�����}T��E�|p�6�I/���~o!L��� Dlma��z/��TOV�����x��~Vs�f^������:�t}^�sٌ�&�4�R���d^!�I4IaX��������٥�0r��NF<5�O9eC~�[�xp7q�c#H2�c|�0+��	6�R��g����%/�\e�y3=�T��%�l�]QԿ�u�]lG��8���גC��~�h*�nIv>��r�^����~EZ�LV�'`X{ �xԂ�g��Pw͹��2���9��`��֒��e��T5�xL�7�qG�i�8o=��@����'�\�~霾(�V��W֩t�k"���^�Ǌ��?w��d��b��Qw����Ik�5��;sUMSVغ16�0\$�Y0�u �?kն)1���r�D�Lٖ)u��2^B� »UX�2��H?dd�s}c-��W��Ww��y�7�x0ɗ�jW��;X�fr�i��tX����Di[�W���|W#q�.���q����E��\LlF���K�S�A��R���!.��x
Ƙ�����`��ڱJ�T��b�p}���f<���,Y䏶\�H�}��VI�`������˫�y��/�C�vZٙ�?:@��W�	/��o^��*��q��=t�eσ��P���ꗒ'��-)Ͷ�p�����ҹ��ͭ�]�@������w�\�آ��'揉C���w�$�BZ��ؠZ��q8�o�r=� �W�Z��/~F!$���r25���:��=���a3|����X�T��L���Vg��Y;O �4�q���(�{]��cIo�������Ge���#�p��x&�� �������Lƨ�>�+rST�Q��	K(�F$W|Iٞ���|A��yn�ԉ���l�ވ�ث)2������w?�Z�ộ�R]k�ʥ*�w�e�HW� A��D0�q3Ub�yZ�^�p���ߨB�@x��a}H����Ǎ�z�g��)�� W�gI��+���`�r���X�� ������+c����/��xy�@��&>(�5F@��ȥ\��^tA�X,vS�@���\o�)�ղ��Uo#娋�5rN��{�-��҆���X0�ѧ֡$�h7-�LgE3^&Hx�$oN���=���ͨ!�9k����k�ܶ_y2���tYxB�y����3�%��-M���xH0j��]O3Y�]�����P�w J�����.r�h�t�˛����a���2�qr�lL��w��C~�ߚ�y���A��#�2I�����]�s��`܇݃b���1�� ��Y������5n�H[��c����/�k�.ȟf�@�<=3���������X!Z2ͩ����P�(����RiX�� ,w��[=�8;Ao0���_r��L�4d:9�7'%\��?����"�3T}h���$/�D�q�FV^�S�������n�QN0�f,�Pp�H����Q�.�c��d��L���bb%�=h �BڽJ�S0|��ɒ4Z��jW?M�Č����s�ՋE��w@Ҕ�d�%��w��aP�*���)3��'>��kV��ؔ�3�6�Au3s_��$�:f=�l΁!�ӯa�e�}�Ij0[Z_K��`Dj��1S]�A+"��-�
��^�~2�k���W�Ij��N�.}��gMڥ�?�&�K��aێ۬��|l�c˾��M��׍�d|K���߄sӆF��O���@h���S�Їx���v�*x)B_[��L������(����8o�H�$��s����s�㉁)��d��Xᚄ�H��<D(R��B��z7��ద]7�>��.A����g�N!:˫����������U�����N����[��Ӕ�s�{��c�7qq�$`��%1w�GD}]R3�G�۽뤊�59����� _q�X��\�1e�Fg�P O%���%�+� j\ЫZ\T˕z�wɒ�xr+1|�cMb�Q)��6�Mh(L���߽.�	(���k�&]k	J� �����[C\�vpO�3j�f �c.9Lz�֯�$_��פ��|ҫF?5^ݮ����Oo��=7���Rڷ�RF�`#�����ŶMa5��~U�27�6������S�($�I)/�z�O[]����~Ȉ]�n����%]�,m�u.lK-B������C=?k�Q>R%|���OȀ�~yk9� ��)n�� z�*f�DX÷��y�C}�k"�_�ͥ9�=���b%�e� �%�0�̳��$N0�E���	��!mu
���.���x
��+�����9&���g���wc�0K/�:X����!�a7)(��k�����x5P(v󩏈�	VZ:\ �B�� η����|(��P���u0���y)�P��ɟ����6��Rf��}գ	��so2�W8�S֨yX��7G��8��yP�¼�f�N    pL=GVf*��p�b�}�/(A*�C5_0��G��X�B �F\�؊x��iǒe��L�#`�Ͳ�� t�w��F��ԛ�IT&p�53�˴V?S���UX�C��Bp;���C\,�T6��Jcb�F8зdy�t��W��>p�����|?�����h?ϧw1j`bpO��X�F�z�-U�N�a�"��T��N�l�$O ��+*q�gXe,������ٯW���М!�*���Z�&p���TV�g��+��ؕR���f{�3��]��@�~գ�� ���������S�6X��7��HgG'���4nHʴJW)��Bkx#[m���eI����s�2�D;��'/�`#E�SE=�)N<��n�6c����>���Z�����y��1��������	!���5���&)x���/��{�NR��R�@��ׁ�˙&ޞ�����n@A���,q�&��D^"^�@+Jf���N�sb��^�R�#5���1�-�ă$�TО��q7�7��h覦j��}�ӿ�Ȇ�j�ǹ��kλ���d�⨖��:L,8��k�^܈-\�{ �1�~R����5���~4uN�I���H��1*\&蜈�5K��wf�5��D��us��ތӤs��,М������/7��&��'��X�L��E��;�>;^оW�Ϭ-�)�&$}7�x�,�2�����cl�t#:�hN��;�`�a[}�O�Ȧ1fk:6��mp�Epǽ4*�����&�<L$6^�%@�OX��� �@��~.WDGŒږQa����zՊZ9^~���|���� �[A�I&���Ί�vV1������^r��������SB$��X�E�Lz*�����`f ����x,����%e	|Vm��f_P��N]搦-NA�\Aq�u����J�#r�ڠ���x�1���8�S��7�1o
4��̡�j���d2�4�-Ơ�Q�q�������,�EX1����v�ƶx�u��ق���A��\�����,l�J�bg���㣜G4DZ�wJ���Z�ޏ�S�N�Ϭύ�(ڒ\��0�z[������"�<#�5��)h���uyc�帡$��8J�T��� 2G8��K�6�䕵kg��͝ߴ��V���IRc�m�7���\��HSK�舊�L���%(�Ec/Y|e�a��������&��;P��Z�n���Y��1�������5&a���/���f�sr��xi�a.��
��v蛋��A��ܧ�Ҡ�/��j�oHb��q\p�4�uU�k."�2%���z��
��|rD+���^�<�j1}����~$e˻�q^����Py�4���{7W㶛�|+j5X�W^��+�|P륕#Ř�3g"E�xh��V;'�&��j�h�������.X/.�;�ɢo@\˷�l��Ҁ�����%�髭(A�c������{��;�J&�&�雛�S�2� r���D�����߄c���b'�c�D�4 ��s���\|��`~z�];���,C�qN�-S֐ ˣ�f�	G'�X^����|n����K�&������ݓl��j���[���������������9�|p�\Z�����"mr!�6D"R
p6��)y�uP��<������P��^����%���I@%��e)��g�#
�< y� <�:�yҡ���'P�4��P՚���J��v�A��n� ���;���(B67�90��~-cRQg���~R���� Aԍ9���j��3nR
�dh��3�Q-]6�D�I�)֚���c�Hnb0���_��B��)e�P�h&��<�E���%_����݊�D�qÈK�B��3ݘ��8͸X
�)ABrZ�+#��f�M�!��%T$�՗X,v{�Rƕ��.�R�2�@tR:��3Ə^�?���"bN`�e2d�րb���cU�6������a��5{���u�2�tlP���
��%{�51%�1,��eb&�iZ����t��Zt'���m� l�0���lu� �����JS�c���,�,�&$��m�Y.��j*��jO�Ahw�����}��2:�G���M7��^�V�E�6h�5<&�)lR5����Ӛ(Q}�-�[�% 5�k��RT�E�q �=Iw����C��$`�#�,srO��dGQ��4�����G@� *���,�k�lߞF��'<�G�h�ʙ��o���+��dǗ���n�#=���➤֖b�;q�� ��Ń.I.s�N�Bp�Qx����8�n�V����)���d��X2x�ⱨ���	�.��
��9��'�ǜ`�y�;�����8��<�Cߠ˃�) ��֙�j=md;��
hҨ@��{��z�wBG�n�����ܧ.{ʬK���6fs�mH�%]U<X]��9Aۡi�gH��	bSW]~	�����G�ݫv{9�

���C���>��M�D)�WA�]�����t��.��;��W�Q�+�Jc��f4 IcҒ��z�aAs�����bɳ�=}Nr�PWD9.m��oq��χ9_��\�)���`� �.	��"�@KR��&o����c���9���+9��4͚�c����;^JK���W
���	��Dܷ�p��&�wkxc�D5�ӌ�7N�E��K�dمD�W�%B���&\�r�j��&3�m����F��#��A��~�xl�6N"tπ#��d`0IKOX��^Z�����uW���GbG<QV��LyՊ�e4�����<	��Ѿ*Wu 1�=���F �E�W���8���X(� H D]G2�ME_�ec �~�F��iE��*y���>�d"��5���3#.���&~;�D�����L0ib>��#�{���5�a9��O/.��Z�)4�0���t9�	@��.b0�'��(��yۋ���:H���@wB�"��\�Q�b	�.�w�P�-����m5�pYqg2�+#"�):�(��_\�ʯ��}���r��_�����=��J+YwV�7Iy��.��O\q�>y��dmY`��k	gÓL���e�������^�WH�OY�(�t�#�Q���8'�=�uO:U� `�4�R�L�=0�B��U�ٓ@(���{�"�����P�\��f�1z4��;;}����^���2��)n���X�,��'	 �j6ƞ"���-��hU֮��ThZH�z@�\'|.;F"Ӌ�d��W��'�؎�Z�w���Սt�X �ވK��)c���`����:ڮ�z������\E�=���>,��C:�(�P��A�$���4�����־w1x�N���W!���bzf�A�JV�A�׉{�uV�܋�;{EGr��V��g��$����5J^R�I��p�F���t���é`V^��,%�k�3��z`8��y.�=�=݊S�[p�ˋ����/��ɫ�.��Fo��N���m�4.��	�����99�Cf{�����TM��_�!�(9ґ��h�5'�����n������<u���іH��o��NQ��U��/����P��P�[g���vIĎѩ���@��)qÙeF�R=2]�/��O땢dH�Y��e6�wZ�!63�=��uf�5 �$.�kt?a]m�ԁ��%�vj����?�e�R���n���9�۵Ndb�O0`��)/�N?lX���y���}�/+�Aq@ͨÆ4w�8��dݜ{���L'�JlĘ��<�7Y����%]M��4>z���X�v���]G!������#x�trX�����vR=��5tf�@²�<%R�\@Y�}&u'�f�v ۦ�b��� �P���'@�3���3���_͏��~w|c"���No��g���7�U�:��h�UTòݠ.=K�Πd�$t/i\�T��m��b֕����NJ˞�ȌA��,43��	�H��˕V��(/���+�q�龑�^/�1��$�]�w��w"���i���eh�K�ҫ�� !���R���G�L1�������4l���SO�S{D�<��O����'�Q�����7���	S��y^^�˕Hd�ͺ�'᳡E|�5 �%˫��[��7�G߀��\��!��=�LOG�b0�$!�\^�$���f�����sY�x�k-��z�?L�Az캝�dO� �i��#��˻��0�bJ�g���,gA�'�a����B�>�/���rXW���ڦ�zd!�孯�H��
��NIv�J��Z�_c>�'aw�Tڋ�s\�ޠ�8T\Rns1�;D�MV=�Œ�欚JW�ҫ�g�����7��E�튅M��K�w��FE��Ģ��PF�t}]����)�s�G�u]���b0�BBB�)D-��*�W�!^�����n����0+�gi,�wX�Oڈ���!(�Do����x�x��~�`�VUsɮ�1&��Lņ�+�m��(�w�Q)���!�_�\�5�����R�p���mh��7������8����<�dI�D�L{�C=�2|�(��2�����O�cd�uq�JO%߄�g��MI:y�H^���,4���g(b=O2����cBO;:�{�,n���>Gvd�� a�dV��c�p?��g-�G�QW�{��҃kD��\��/�ص�mԌ�튦���+1-�n����UA٩����3�1�2bQ���E֘���K��@w������ۓqY��8�3̆N^�H�<��WW���%e|��$�w���{"�e7�]�����U��I�7�z�n�-�be�����̮(-�|�4s-�6�`�UB��AK;'�ƃg�tj(>!�W�a\��|+���;}�b뷚[�!>v졢�����w9��t�����i\��J���3�F"0�l=�5�UD��N?��(۲��t�38$������bfoբ0�׿:�;|�'k7���'�/3��\Y���B�w�O�jw��#�9�/����V|E Y��	�;�v.�z~"�q�+!Зl��'Q�?{�m��PV����\�8l�}E��t�$?V�Ib/TF�I���[�;��3'|Y��|�)T�%�2X+D��B��/��������C~<*_��(��������?[]�5c蛋���al���~�e��,_2�=�&�Wf��lz�[�sҬ)���㛃@TU�����mt�U�Ǯe*u�g@��#�5a��)����v���_�U-����<�|խ����1���-J�O�u�����u���`�n�a���u�B�U�"�Dx�G���\���=縷l��� �"�w������2D�(T]���w�%&�������-N�c�����Y7�d�<�m>q�ě��x�|����_��qp���i^E�cr�Rz�5h�삙sN���^�|-j����~i���Bc��E����{s�)��JPw�|�>�&P�p��Q6���!�$c�f�/���ú��k+�Y'A?IC!.3�&�]�u��͏L^HT���
ĸ��E2r�S���@�k0���vG@�Rwb�SFD�smg��~��;p���@�=(3��Jw�o:U��rE��ڎM�@@%�w�zkBC��6G�$Y����0|�lt�����R�eLY�z�阧m��Q�l�����>}��cV��$�:a�]/�'f��5����%���~V�m���	��G��������. �z�j��N��"2���c�+��/يpT�Y$L22����_���"�:�W��k�ӠO���5�b�i�����fxV]��s���r���Qr���������-�x���6��M��s�����gr�]z�C���P�4���Bc�CGoQh�/�a@H�r�N�i��;�$�lA!��MM]JA{�r�!d����)�ZU�I*�a��dE���rQ_�jgk�}Z�LI�8<s6��G
�B�k��W��YʜV��|Ep���h}ϊߟ\�����z��C�{<�˰4jz���K[M�H5��2堢򸢴(CXr�'я�TԂk�T��cp7���%�&�1$�R��,��+�O@�7�y$�/�9�̼��Z|,���<4hU���~([{͟�e�K��GB"�h�`�����N�<M�rHn\��t$���@�d�3���wa^5�f!�D�9�/�C9e
Rei���~	C<��Ig�d��7��8ʘ�h&��iF�3x,�� 7(��n79� z�:�����*��i�ݷ���������O�E���@��!r�)/�G�ڔ��A�A}7�����k�5� =�a�X���fU��Q�ܻ�^"!�)�=��+e�w�/xH���3��:4"��zn^��@��ԈO�&��۽u�l�ܨmң�w�[��X���D��Ҙ�Z�zV�%4��/�~�
���5�ۧD��0�uiOo�����͝pۼٹ�W�4B�s��'J�����.�"��Uz�|����R�M��E�T*�_�۞/G��P�� �p���y��ӂG��.|9�k;%������Kt���ĕe	ǅv����!DC����A&�K	<>h=/,a F�bW�V��b�ta�M攂�6�ϫ�4Ԟ�'1R�/�0$3���%�B������ nteoQ�2������?)�y��Տ9"�,�q���d$�@��£D߫���2?}{���+���N�3�[U���V?� �������AS7��vu�`������_?̎/˔]L(�Xd_"ǯK��ܯ�P���%-tD�+�\�CB��ޙ���K�d�E��E �L�� ��նY�q�	[e%�M��K���1j}y$$0��W3y^u�;\S6M�����Ó+[݉�6F��A��%�軵��ͥ�\~�J��[�4�����;a���*���3����Ao|`�R��,�Q '��dȾQ@���G���\R(�ƠL�����X��R�7^�a	�3�"��P5[�\M�X�����K�g�yA<���"&;�w�U����w�R[W��sSWa��pHr4����'a�Ѳ�1�S*'�W���f+�c	����e��>��Z�V��I��9��������������]#'�Z�Ć���+F-9��Ѩ+a}��0�q ˝ę�����"�߯v�;}����DK��N���5���W]e��T��,��މvv�!���w�'o���_�*�З�(\7]`5��\y)9M"����ew݂�r��,�g�H|�G��M�hB�}�2�IM����xun�(�_	���P>H.���@�����T��۞�X#4�q�KNـ�-CI�����r|M�0�q �b�����+ZQR�������IJγmp>Nt��-���8�y�r�myz}@��Q����	dƅ!%�U� �pC��P�bø�y]�=��`�h,p�1���jC��	�a����v�dI��}����+WL\1���̃PH��`k�J�è��|��$��߁���,�8�㺡#fRi6��[�����gަ�0d��_�;&ހٹ��K��eS2γ�<;6�������
r��4����=�pVO�ąO��S.=f	�8c¶H�D��Mq�$W���mS��tA��ɬ�<k�˲HcꚇD�^*��"�����e��&�N��e�uS�i��Э8
��u.��d$�^��Ib��ĵ�c4�9*���bV�;&��I��OĝX��	�����޹֩����J��G8�uS<Q��;�.P������2�p�_?��8¦;J���tY'!/6'2��?3��jR��r�6���ބ�x�ǣS�^^��;���[4�Q(�7��c#݂]�v��l�D�=	�ͬ^D���םj޻���G�R+�����,aLm�/�̅q��$�E��%Y��9(Վ�"\2.}�y�x>��b�u�Jp<���%�^�rD
S �(�djh��7K*�݇�Xx �X�^���Y���� �]T%��S���(�^�j>1ugƦ#L��Ա����~�1�+����^���h�y�`1��1dܻ*��[��eN�b)�#�4"�~�C'�;k��2[w���
J�U���ŉ":� G:j_��r��ܹ#[4��a�.��]b�i�rt�y�.��DuB�B�[v��.���q���zd�]�t�@�n.�1˛#��5aR.h#�&�l��'��CI��,h�g����ؑ���1B�;?M����.��MP?���t���P+���B2�ႶZ
0��T�X�	��MDA^D%0��&�K�҄a�� ����^�?X��Ún����I!(N�pC5�B�]Δ����?X�;�CAW�3k���u�,~�W�RWX Q�L�8�Էo�;UC�hPҎ��e;<_]ފ������l[U��s�A�W2L�ӧ�g(�r�&�u?*@0�+Xq�
۵��/h���ߖ� ����yEy�Ћ��M�{�,z)1� ��i�]�U���ʥ^O����Y�Ӈ��J�s�rs�2��Vy%J~��#�z��lj�EN���FȂ*Σ�B���ώдI�R�l�?�G
ق>E�����=��@���N��K����G>�N�"C��'{� �]�!3�C2��_/|�C&2�W��x�y�#���.�S	�Zc�V�Uw띬�A���HZN�h�W�F�p��X�[��lo!�q.��LT�$(H�¦�P�O=�ש4�0����M/��Zw��>dQ�~�8m������lgT�9�����:��� M�*&��W�$p�-���